-- megafunction wizard: %LPM_MUX%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: lpm_mux 

-- ============================================================
-- File Name: lpm_muxVDM.vhd
-- Megafunction Name(s):
-- 			lpm_mux
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 9.1 Build 222 10/21/2009 SJ Web Edition
-- ************************************************************


--Copyright (C) 1991-2009 Altera Corporation
--Your use of Altera Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Altera Program License 
--Subscription Agreement, Altera MegaCore Function License 
--Agreement, or other applicable license agreement, including, 
--without limitation, that your use is for the sole purpose of 
--programming logic devices manufactured by Altera and sold by 
--Altera or its authorized distributors.  Please refer to the 
--applicable agreement for further details.


LIBRARY ieee;
USE ieee.std_logic_1164.all;

LIBRARY lpm;
USE lpm.lpm_components.all;

ENTITY lpm_muxVDM IS
	PORT
	(
		data0x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data10x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data11x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data12x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data13x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data14x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data15x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data1x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data2x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data3x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data4x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data5x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data6x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data7x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data8x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		data9x		: IN STD_LOGIC_VECTOR (127 DOWNTO 0);
		sel		: IN STD_LOGIC_VECTOR (3 DOWNTO 0);
		result		: OUT STD_LOGIC_VECTOR (127 DOWNTO 0)
	);
END lpm_muxVDM;


ARCHITECTURE SYN OF lpm_muxvdm IS

--	type STD_LOGIC_2D is array (NATURAL RANGE <>, NATURAL RANGE <>) of STD_LOGIC;

	SIGNAL sub_wire0	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire2	: STD_LOGIC_2D (15 DOWNTO 0, 127 DOWNTO 0);
	SIGNAL sub_wire3	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire4	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire5	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire6	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire7	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire8	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire9	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire10	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire11	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire12	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire13	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire14	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire15	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire16	: STD_LOGIC_VECTOR (127 DOWNTO 0);
	SIGNAL sub_wire17	: STD_LOGIC_VECTOR (127 DOWNTO 0);

BEGIN
	sub_wire17    <= data0x(127 DOWNTO 0);
	sub_wire16    <= data1x(127 DOWNTO 0);
	sub_wire15    <= data2x(127 DOWNTO 0);
	sub_wire14    <= data3x(127 DOWNTO 0);
	sub_wire13    <= data4x(127 DOWNTO 0);
	sub_wire12    <= data5x(127 DOWNTO 0);
	sub_wire11    <= data6x(127 DOWNTO 0);
	sub_wire10    <= data7x(127 DOWNTO 0);
	sub_wire9    <= data8x(127 DOWNTO 0);
	sub_wire8    <= data9x(127 DOWNTO 0);
	sub_wire7    <= data10x(127 DOWNTO 0);
	sub_wire6    <= data11x(127 DOWNTO 0);
	sub_wire5    <= data12x(127 DOWNTO 0);
	sub_wire4    <= data13x(127 DOWNTO 0);
	sub_wire3    <= data14x(127 DOWNTO 0);
	result    <= sub_wire0(127 DOWNTO 0);
	sub_wire1    <= data15x(127 DOWNTO 0);
	sub_wire2(15, 0)    <= sub_wire1(0);
	sub_wire2(15, 1)    <= sub_wire1(1);
	sub_wire2(15, 2)    <= sub_wire1(2);
	sub_wire2(15, 3)    <= sub_wire1(3);
	sub_wire2(15, 4)    <= sub_wire1(4);
	sub_wire2(15, 5)    <= sub_wire1(5);
	sub_wire2(15, 6)    <= sub_wire1(6);
	sub_wire2(15, 7)    <= sub_wire1(7);
	sub_wire2(15, 8)    <= sub_wire1(8);
	sub_wire2(15, 9)    <= sub_wire1(9);
	sub_wire2(15, 10)    <= sub_wire1(10);
	sub_wire2(15, 11)    <= sub_wire1(11);
	sub_wire2(15, 12)    <= sub_wire1(12);
	sub_wire2(15, 13)    <= sub_wire1(13);
	sub_wire2(15, 14)    <= sub_wire1(14);
	sub_wire2(15, 15)    <= sub_wire1(15);
	sub_wire2(15, 16)    <= sub_wire1(16);
	sub_wire2(15, 17)    <= sub_wire1(17);
	sub_wire2(15, 18)    <= sub_wire1(18);
	sub_wire2(15, 19)    <= sub_wire1(19);
	sub_wire2(15, 20)    <= sub_wire1(20);
	sub_wire2(15, 21)    <= sub_wire1(21);
	sub_wire2(15, 22)    <= sub_wire1(22);
	sub_wire2(15, 23)    <= sub_wire1(23);
	sub_wire2(15, 24)    <= sub_wire1(24);
	sub_wire2(15, 25)    <= sub_wire1(25);
	sub_wire2(15, 26)    <= sub_wire1(26);
	sub_wire2(15, 27)    <= sub_wire1(27);
	sub_wire2(15, 28)    <= sub_wire1(28);
	sub_wire2(15, 29)    <= sub_wire1(29);
	sub_wire2(15, 30)    <= sub_wire1(30);
	sub_wire2(15, 31)    <= sub_wire1(31);
	sub_wire2(15, 32)    <= sub_wire1(32);
	sub_wire2(15, 33)    <= sub_wire1(33);
	sub_wire2(15, 34)    <= sub_wire1(34);
	sub_wire2(15, 35)    <= sub_wire1(35);
	sub_wire2(15, 36)    <= sub_wire1(36);
	sub_wire2(15, 37)    <= sub_wire1(37);
	sub_wire2(15, 38)    <= sub_wire1(38);
	sub_wire2(15, 39)    <= sub_wire1(39);
	sub_wire2(15, 40)    <= sub_wire1(40);
	sub_wire2(15, 41)    <= sub_wire1(41);
	sub_wire2(15, 42)    <= sub_wire1(42);
	sub_wire2(15, 43)    <= sub_wire1(43);
	sub_wire2(15, 44)    <= sub_wire1(44);
	sub_wire2(15, 45)    <= sub_wire1(45);
	sub_wire2(15, 46)    <= sub_wire1(46);
	sub_wire2(15, 47)    <= sub_wire1(47);
	sub_wire2(15, 48)    <= sub_wire1(48);
	sub_wire2(15, 49)    <= sub_wire1(49);
	sub_wire2(15, 50)    <= sub_wire1(50);
	sub_wire2(15, 51)    <= sub_wire1(51);
	sub_wire2(15, 52)    <= sub_wire1(52);
	sub_wire2(15, 53)    <= sub_wire1(53);
	sub_wire2(15, 54)    <= sub_wire1(54);
	sub_wire2(15, 55)    <= sub_wire1(55);
	sub_wire2(15, 56)    <= sub_wire1(56);
	sub_wire2(15, 57)    <= sub_wire1(57);
	sub_wire2(15, 58)    <= sub_wire1(58);
	sub_wire2(15, 59)    <= sub_wire1(59);
	sub_wire2(15, 60)    <= sub_wire1(60);
	sub_wire2(15, 61)    <= sub_wire1(61);
	sub_wire2(15, 62)    <= sub_wire1(62);
	sub_wire2(15, 63)    <= sub_wire1(63);
	sub_wire2(15, 64)    <= sub_wire1(64);
	sub_wire2(15, 65)    <= sub_wire1(65);
	sub_wire2(15, 66)    <= sub_wire1(66);
	sub_wire2(15, 67)    <= sub_wire1(67);
	sub_wire2(15, 68)    <= sub_wire1(68);
	sub_wire2(15, 69)    <= sub_wire1(69);
	sub_wire2(15, 70)    <= sub_wire1(70);
	sub_wire2(15, 71)    <= sub_wire1(71);
	sub_wire2(15, 72)    <= sub_wire1(72);
	sub_wire2(15, 73)    <= sub_wire1(73);
	sub_wire2(15, 74)    <= sub_wire1(74);
	sub_wire2(15, 75)    <= sub_wire1(75);
	sub_wire2(15, 76)    <= sub_wire1(76);
	sub_wire2(15, 77)    <= sub_wire1(77);
	sub_wire2(15, 78)    <= sub_wire1(78);
	sub_wire2(15, 79)    <= sub_wire1(79);
	sub_wire2(15, 80)    <= sub_wire1(80);
	sub_wire2(15, 81)    <= sub_wire1(81);
	sub_wire2(15, 82)    <= sub_wire1(82);
	sub_wire2(15, 83)    <= sub_wire1(83);
	sub_wire2(15, 84)    <= sub_wire1(84);
	sub_wire2(15, 85)    <= sub_wire1(85);
	sub_wire2(15, 86)    <= sub_wire1(86);
	sub_wire2(15, 87)    <= sub_wire1(87);
	sub_wire2(15, 88)    <= sub_wire1(88);
	sub_wire2(15, 89)    <= sub_wire1(89);
	sub_wire2(15, 90)    <= sub_wire1(90);
	sub_wire2(15, 91)    <= sub_wire1(91);
	sub_wire2(15, 92)    <= sub_wire1(92);
	sub_wire2(15, 93)    <= sub_wire1(93);
	sub_wire2(15, 94)    <= sub_wire1(94);
	sub_wire2(15, 95)    <= sub_wire1(95);
	sub_wire2(15, 96)    <= sub_wire1(96);
	sub_wire2(15, 97)    <= sub_wire1(97);
	sub_wire2(15, 98)    <= sub_wire1(98);
	sub_wire2(15, 99)    <= sub_wire1(99);
	sub_wire2(15, 100)    <= sub_wire1(100);
	sub_wire2(15, 101)    <= sub_wire1(101);
	sub_wire2(15, 102)    <= sub_wire1(102);
	sub_wire2(15, 103)    <= sub_wire1(103);
	sub_wire2(15, 104)    <= sub_wire1(104);
	sub_wire2(15, 105)    <= sub_wire1(105);
	sub_wire2(15, 106)    <= sub_wire1(106);
	sub_wire2(15, 107)    <= sub_wire1(107);
	sub_wire2(15, 108)    <= sub_wire1(108);
	sub_wire2(15, 109)    <= sub_wire1(109);
	sub_wire2(15, 110)    <= sub_wire1(110);
	sub_wire2(15, 111)    <= sub_wire1(111);
	sub_wire2(15, 112)    <= sub_wire1(112);
	sub_wire2(15, 113)    <= sub_wire1(113);
	sub_wire2(15, 114)    <= sub_wire1(114);
	sub_wire2(15, 115)    <= sub_wire1(115);
	sub_wire2(15, 116)    <= sub_wire1(116);
	sub_wire2(15, 117)    <= sub_wire1(117);
	sub_wire2(15, 118)    <= sub_wire1(118);
	sub_wire2(15, 119)    <= sub_wire1(119);
	sub_wire2(15, 120)    <= sub_wire1(120);
	sub_wire2(15, 121)    <= sub_wire1(121);
	sub_wire2(15, 122)    <= sub_wire1(122);
	sub_wire2(15, 123)    <= sub_wire1(123);
	sub_wire2(15, 124)    <= sub_wire1(124);
	sub_wire2(15, 125)    <= sub_wire1(125);
	sub_wire2(15, 126)    <= sub_wire1(126);
	sub_wire2(15, 127)    <= sub_wire1(127);
	sub_wire2(14, 0)    <= sub_wire3(0);
	sub_wire2(14, 1)    <= sub_wire3(1);
	sub_wire2(14, 2)    <= sub_wire3(2);
	sub_wire2(14, 3)    <= sub_wire3(3);
	sub_wire2(14, 4)    <= sub_wire3(4);
	sub_wire2(14, 5)    <= sub_wire3(5);
	sub_wire2(14, 6)    <= sub_wire3(6);
	sub_wire2(14, 7)    <= sub_wire3(7);
	sub_wire2(14, 8)    <= sub_wire3(8);
	sub_wire2(14, 9)    <= sub_wire3(9);
	sub_wire2(14, 10)    <= sub_wire3(10);
	sub_wire2(14, 11)    <= sub_wire3(11);
	sub_wire2(14, 12)    <= sub_wire3(12);
	sub_wire2(14, 13)    <= sub_wire3(13);
	sub_wire2(14, 14)    <= sub_wire3(14);
	sub_wire2(14, 15)    <= sub_wire3(15);
	sub_wire2(14, 16)    <= sub_wire3(16);
	sub_wire2(14, 17)    <= sub_wire3(17);
	sub_wire2(14, 18)    <= sub_wire3(18);
	sub_wire2(14, 19)    <= sub_wire3(19);
	sub_wire2(14, 20)    <= sub_wire3(20);
	sub_wire2(14, 21)    <= sub_wire3(21);
	sub_wire2(14, 22)    <= sub_wire3(22);
	sub_wire2(14, 23)    <= sub_wire3(23);
	sub_wire2(14, 24)    <= sub_wire3(24);
	sub_wire2(14, 25)    <= sub_wire3(25);
	sub_wire2(14, 26)    <= sub_wire3(26);
	sub_wire2(14, 27)    <= sub_wire3(27);
	sub_wire2(14, 28)    <= sub_wire3(28);
	sub_wire2(14, 29)    <= sub_wire3(29);
	sub_wire2(14, 30)    <= sub_wire3(30);
	sub_wire2(14, 31)    <= sub_wire3(31);
	sub_wire2(14, 32)    <= sub_wire3(32);
	sub_wire2(14, 33)    <= sub_wire3(33);
	sub_wire2(14, 34)    <= sub_wire3(34);
	sub_wire2(14, 35)    <= sub_wire3(35);
	sub_wire2(14, 36)    <= sub_wire3(36);
	sub_wire2(14, 37)    <= sub_wire3(37);
	sub_wire2(14, 38)    <= sub_wire3(38);
	sub_wire2(14, 39)    <= sub_wire3(39);
	sub_wire2(14, 40)    <= sub_wire3(40);
	sub_wire2(14, 41)    <= sub_wire3(41);
	sub_wire2(14, 42)    <= sub_wire3(42);
	sub_wire2(14, 43)    <= sub_wire3(43);
	sub_wire2(14, 44)    <= sub_wire3(44);
	sub_wire2(14, 45)    <= sub_wire3(45);
	sub_wire2(14, 46)    <= sub_wire3(46);
	sub_wire2(14, 47)    <= sub_wire3(47);
	sub_wire2(14, 48)    <= sub_wire3(48);
	sub_wire2(14, 49)    <= sub_wire3(49);
	sub_wire2(14, 50)    <= sub_wire3(50);
	sub_wire2(14, 51)    <= sub_wire3(51);
	sub_wire2(14, 52)    <= sub_wire3(52);
	sub_wire2(14, 53)    <= sub_wire3(53);
	sub_wire2(14, 54)    <= sub_wire3(54);
	sub_wire2(14, 55)    <= sub_wire3(55);
	sub_wire2(14, 56)    <= sub_wire3(56);
	sub_wire2(14, 57)    <= sub_wire3(57);
	sub_wire2(14, 58)    <= sub_wire3(58);
	sub_wire2(14, 59)    <= sub_wire3(59);
	sub_wire2(14, 60)    <= sub_wire3(60);
	sub_wire2(14, 61)    <= sub_wire3(61);
	sub_wire2(14, 62)    <= sub_wire3(62);
	sub_wire2(14, 63)    <= sub_wire3(63);
	sub_wire2(14, 64)    <= sub_wire3(64);
	sub_wire2(14, 65)    <= sub_wire3(65);
	sub_wire2(14, 66)    <= sub_wire3(66);
	sub_wire2(14, 67)    <= sub_wire3(67);
	sub_wire2(14, 68)    <= sub_wire3(68);
	sub_wire2(14, 69)    <= sub_wire3(69);
	sub_wire2(14, 70)    <= sub_wire3(70);
	sub_wire2(14, 71)    <= sub_wire3(71);
	sub_wire2(14, 72)    <= sub_wire3(72);
	sub_wire2(14, 73)    <= sub_wire3(73);
	sub_wire2(14, 74)    <= sub_wire3(74);
	sub_wire2(14, 75)    <= sub_wire3(75);
	sub_wire2(14, 76)    <= sub_wire3(76);
	sub_wire2(14, 77)    <= sub_wire3(77);
	sub_wire2(14, 78)    <= sub_wire3(78);
	sub_wire2(14, 79)    <= sub_wire3(79);
	sub_wire2(14, 80)    <= sub_wire3(80);
	sub_wire2(14, 81)    <= sub_wire3(81);
	sub_wire2(14, 82)    <= sub_wire3(82);
	sub_wire2(14, 83)    <= sub_wire3(83);
	sub_wire2(14, 84)    <= sub_wire3(84);
	sub_wire2(14, 85)    <= sub_wire3(85);
	sub_wire2(14, 86)    <= sub_wire3(86);
	sub_wire2(14, 87)    <= sub_wire3(87);
	sub_wire2(14, 88)    <= sub_wire3(88);
	sub_wire2(14, 89)    <= sub_wire3(89);
	sub_wire2(14, 90)    <= sub_wire3(90);
	sub_wire2(14, 91)    <= sub_wire3(91);
	sub_wire2(14, 92)    <= sub_wire3(92);
	sub_wire2(14, 93)    <= sub_wire3(93);
	sub_wire2(14, 94)    <= sub_wire3(94);
	sub_wire2(14, 95)    <= sub_wire3(95);
	sub_wire2(14, 96)    <= sub_wire3(96);
	sub_wire2(14, 97)    <= sub_wire3(97);
	sub_wire2(14, 98)    <= sub_wire3(98);
	sub_wire2(14, 99)    <= sub_wire3(99);
	sub_wire2(14, 100)    <= sub_wire3(100);
	sub_wire2(14, 101)    <= sub_wire3(101);
	sub_wire2(14, 102)    <= sub_wire3(102);
	sub_wire2(14, 103)    <= sub_wire3(103);
	sub_wire2(14, 104)    <= sub_wire3(104);
	sub_wire2(14, 105)    <= sub_wire3(105);
	sub_wire2(14, 106)    <= sub_wire3(106);
	sub_wire2(14, 107)    <= sub_wire3(107);
	sub_wire2(14, 108)    <= sub_wire3(108);
	sub_wire2(14, 109)    <= sub_wire3(109);
	sub_wire2(14, 110)    <= sub_wire3(110);
	sub_wire2(14, 111)    <= sub_wire3(111);
	sub_wire2(14, 112)    <= sub_wire3(112);
	sub_wire2(14, 113)    <= sub_wire3(113);
	sub_wire2(14, 114)    <= sub_wire3(114);
	sub_wire2(14, 115)    <= sub_wire3(115);
	sub_wire2(14, 116)    <= sub_wire3(116);
	sub_wire2(14, 117)    <= sub_wire3(117);
	sub_wire2(14, 118)    <= sub_wire3(118);
	sub_wire2(14, 119)    <= sub_wire3(119);
	sub_wire2(14, 120)    <= sub_wire3(120);
	sub_wire2(14, 121)    <= sub_wire3(121);
	sub_wire2(14, 122)    <= sub_wire3(122);
	sub_wire2(14, 123)    <= sub_wire3(123);
	sub_wire2(14, 124)    <= sub_wire3(124);
	sub_wire2(14, 125)    <= sub_wire3(125);
	sub_wire2(14, 126)    <= sub_wire3(126);
	sub_wire2(14, 127)    <= sub_wire3(127);
	sub_wire2(13, 0)    <= sub_wire4(0);
	sub_wire2(13, 1)    <= sub_wire4(1);
	sub_wire2(13, 2)    <= sub_wire4(2);
	sub_wire2(13, 3)    <= sub_wire4(3);
	sub_wire2(13, 4)    <= sub_wire4(4);
	sub_wire2(13, 5)    <= sub_wire4(5);
	sub_wire2(13, 6)    <= sub_wire4(6);
	sub_wire2(13, 7)    <= sub_wire4(7);
	sub_wire2(13, 8)    <= sub_wire4(8);
	sub_wire2(13, 9)    <= sub_wire4(9);
	sub_wire2(13, 10)    <= sub_wire4(10);
	sub_wire2(13, 11)    <= sub_wire4(11);
	sub_wire2(13, 12)    <= sub_wire4(12);
	sub_wire2(13, 13)    <= sub_wire4(13);
	sub_wire2(13, 14)    <= sub_wire4(14);
	sub_wire2(13, 15)    <= sub_wire4(15);
	sub_wire2(13, 16)    <= sub_wire4(16);
	sub_wire2(13, 17)    <= sub_wire4(17);
	sub_wire2(13, 18)    <= sub_wire4(18);
	sub_wire2(13, 19)    <= sub_wire4(19);
	sub_wire2(13, 20)    <= sub_wire4(20);
	sub_wire2(13, 21)    <= sub_wire4(21);
	sub_wire2(13, 22)    <= sub_wire4(22);
	sub_wire2(13, 23)    <= sub_wire4(23);
	sub_wire2(13, 24)    <= sub_wire4(24);
	sub_wire2(13, 25)    <= sub_wire4(25);
	sub_wire2(13, 26)    <= sub_wire4(26);
	sub_wire2(13, 27)    <= sub_wire4(27);
	sub_wire2(13, 28)    <= sub_wire4(28);
	sub_wire2(13, 29)    <= sub_wire4(29);
	sub_wire2(13, 30)    <= sub_wire4(30);
	sub_wire2(13, 31)    <= sub_wire4(31);
	sub_wire2(13, 32)    <= sub_wire4(32);
	sub_wire2(13, 33)    <= sub_wire4(33);
	sub_wire2(13, 34)    <= sub_wire4(34);
	sub_wire2(13, 35)    <= sub_wire4(35);
	sub_wire2(13, 36)    <= sub_wire4(36);
	sub_wire2(13, 37)    <= sub_wire4(37);
	sub_wire2(13, 38)    <= sub_wire4(38);
	sub_wire2(13, 39)    <= sub_wire4(39);
	sub_wire2(13, 40)    <= sub_wire4(40);
	sub_wire2(13, 41)    <= sub_wire4(41);
	sub_wire2(13, 42)    <= sub_wire4(42);
	sub_wire2(13, 43)    <= sub_wire4(43);
	sub_wire2(13, 44)    <= sub_wire4(44);
	sub_wire2(13, 45)    <= sub_wire4(45);
	sub_wire2(13, 46)    <= sub_wire4(46);
	sub_wire2(13, 47)    <= sub_wire4(47);
	sub_wire2(13, 48)    <= sub_wire4(48);
	sub_wire2(13, 49)    <= sub_wire4(49);
	sub_wire2(13, 50)    <= sub_wire4(50);
	sub_wire2(13, 51)    <= sub_wire4(51);
	sub_wire2(13, 52)    <= sub_wire4(52);
	sub_wire2(13, 53)    <= sub_wire4(53);
	sub_wire2(13, 54)    <= sub_wire4(54);
	sub_wire2(13, 55)    <= sub_wire4(55);
	sub_wire2(13, 56)    <= sub_wire4(56);
	sub_wire2(13, 57)    <= sub_wire4(57);
	sub_wire2(13, 58)    <= sub_wire4(58);
	sub_wire2(13, 59)    <= sub_wire4(59);
	sub_wire2(13, 60)    <= sub_wire4(60);
	sub_wire2(13, 61)    <= sub_wire4(61);
	sub_wire2(13, 62)    <= sub_wire4(62);
	sub_wire2(13, 63)    <= sub_wire4(63);
	sub_wire2(13, 64)    <= sub_wire4(64);
	sub_wire2(13, 65)    <= sub_wire4(65);
	sub_wire2(13, 66)    <= sub_wire4(66);
	sub_wire2(13, 67)    <= sub_wire4(67);
	sub_wire2(13, 68)    <= sub_wire4(68);
	sub_wire2(13, 69)    <= sub_wire4(69);
	sub_wire2(13, 70)    <= sub_wire4(70);
	sub_wire2(13, 71)    <= sub_wire4(71);
	sub_wire2(13, 72)    <= sub_wire4(72);
	sub_wire2(13, 73)    <= sub_wire4(73);
	sub_wire2(13, 74)    <= sub_wire4(74);
	sub_wire2(13, 75)    <= sub_wire4(75);
	sub_wire2(13, 76)    <= sub_wire4(76);
	sub_wire2(13, 77)    <= sub_wire4(77);
	sub_wire2(13, 78)    <= sub_wire4(78);
	sub_wire2(13, 79)    <= sub_wire4(79);
	sub_wire2(13, 80)    <= sub_wire4(80);
	sub_wire2(13, 81)    <= sub_wire4(81);
	sub_wire2(13, 82)    <= sub_wire4(82);
	sub_wire2(13, 83)    <= sub_wire4(83);
	sub_wire2(13, 84)    <= sub_wire4(84);
	sub_wire2(13, 85)    <= sub_wire4(85);
	sub_wire2(13, 86)    <= sub_wire4(86);
	sub_wire2(13, 87)    <= sub_wire4(87);
	sub_wire2(13, 88)    <= sub_wire4(88);
	sub_wire2(13, 89)    <= sub_wire4(89);
	sub_wire2(13, 90)    <= sub_wire4(90);
	sub_wire2(13, 91)    <= sub_wire4(91);
	sub_wire2(13, 92)    <= sub_wire4(92);
	sub_wire2(13, 93)    <= sub_wire4(93);
	sub_wire2(13, 94)    <= sub_wire4(94);
	sub_wire2(13, 95)    <= sub_wire4(95);
	sub_wire2(13, 96)    <= sub_wire4(96);
	sub_wire2(13, 97)    <= sub_wire4(97);
	sub_wire2(13, 98)    <= sub_wire4(98);
	sub_wire2(13, 99)    <= sub_wire4(99);
	sub_wire2(13, 100)    <= sub_wire4(100);
	sub_wire2(13, 101)    <= sub_wire4(101);
	sub_wire2(13, 102)    <= sub_wire4(102);
	sub_wire2(13, 103)    <= sub_wire4(103);
	sub_wire2(13, 104)    <= sub_wire4(104);
	sub_wire2(13, 105)    <= sub_wire4(105);
	sub_wire2(13, 106)    <= sub_wire4(106);
	sub_wire2(13, 107)    <= sub_wire4(107);
	sub_wire2(13, 108)    <= sub_wire4(108);
	sub_wire2(13, 109)    <= sub_wire4(109);
	sub_wire2(13, 110)    <= sub_wire4(110);
	sub_wire2(13, 111)    <= sub_wire4(111);
	sub_wire2(13, 112)    <= sub_wire4(112);
	sub_wire2(13, 113)    <= sub_wire4(113);
	sub_wire2(13, 114)    <= sub_wire4(114);
	sub_wire2(13, 115)    <= sub_wire4(115);
	sub_wire2(13, 116)    <= sub_wire4(116);
	sub_wire2(13, 117)    <= sub_wire4(117);
	sub_wire2(13, 118)    <= sub_wire4(118);
	sub_wire2(13, 119)    <= sub_wire4(119);
	sub_wire2(13, 120)    <= sub_wire4(120);
	sub_wire2(13, 121)    <= sub_wire4(121);
	sub_wire2(13, 122)    <= sub_wire4(122);
	sub_wire2(13, 123)    <= sub_wire4(123);
	sub_wire2(13, 124)    <= sub_wire4(124);
	sub_wire2(13, 125)    <= sub_wire4(125);
	sub_wire2(13, 126)    <= sub_wire4(126);
	sub_wire2(13, 127)    <= sub_wire4(127);
	sub_wire2(12, 0)    <= sub_wire5(0);
	sub_wire2(12, 1)    <= sub_wire5(1);
	sub_wire2(12, 2)    <= sub_wire5(2);
	sub_wire2(12, 3)    <= sub_wire5(3);
	sub_wire2(12, 4)    <= sub_wire5(4);
	sub_wire2(12, 5)    <= sub_wire5(5);
	sub_wire2(12, 6)    <= sub_wire5(6);
	sub_wire2(12, 7)    <= sub_wire5(7);
	sub_wire2(12, 8)    <= sub_wire5(8);
	sub_wire2(12, 9)    <= sub_wire5(9);
	sub_wire2(12, 10)    <= sub_wire5(10);
	sub_wire2(12, 11)    <= sub_wire5(11);
	sub_wire2(12, 12)    <= sub_wire5(12);
	sub_wire2(12, 13)    <= sub_wire5(13);
	sub_wire2(12, 14)    <= sub_wire5(14);
	sub_wire2(12, 15)    <= sub_wire5(15);
	sub_wire2(12, 16)    <= sub_wire5(16);
	sub_wire2(12, 17)    <= sub_wire5(17);
	sub_wire2(12, 18)    <= sub_wire5(18);
	sub_wire2(12, 19)    <= sub_wire5(19);
	sub_wire2(12, 20)    <= sub_wire5(20);
	sub_wire2(12, 21)    <= sub_wire5(21);
	sub_wire2(12, 22)    <= sub_wire5(22);
	sub_wire2(12, 23)    <= sub_wire5(23);
	sub_wire2(12, 24)    <= sub_wire5(24);
	sub_wire2(12, 25)    <= sub_wire5(25);
	sub_wire2(12, 26)    <= sub_wire5(26);
	sub_wire2(12, 27)    <= sub_wire5(27);
	sub_wire2(12, 28)    <= sub_wire5(28);
	sub_wire2(12, 29)    <= sub_wire5(29);
	sub_wire2(12, 30)    <= sub_wire5(30);
	sub_wire2(12, 31)    <= sub_wire5(31);
	sub_wire2(12, 32)    <= sub_wire5(32);
	sub_wire2(12, 33)    <= sub_wire5(33);
	sub_wire2(12, 34)    <= sub_wire5(34);
	sub_wire2(12, 35)    <= sub_wire5(35);
	sub_wire2(12, 36)    <= sub_wire5(36);
	sub_wire2(12, 37)    <= sub_wire5(37);
	sub_wire2(12, 38)    <= sub_wire5(38);
	sub_wire2(12, 39)    <= sub_wire5(39);
	sub_wire2(12, 40)    <= sub_wire5(40);
	sub_wire2(12, 41)    <= sub_wire5(41);
	sub_wire2(12, 42)    <= sub_wire5(42);
	sub_wire2(12, 43)    <= sub_wire5(43);
	sub_wire2(12, 44)    <= sub_wire5(44);
	sub_wire2(12, 45)    <= sub_wire5(45);
	sub_wire2(12, 46)    <= sub_wire5(46);
	sub_wire2(12, 47)    <= sub_wire5(47);
	sub_wire2(12, 48)    <= sub_wire5(48);
	sub_wire2(12, 49)    <= sub_wire5(49);
	sub_wire2(12, 50)    <= sub_wire5(50);
	sub_wire2(12, 51)    <= sub_wire5(51);
	sub_wire2(12, 52)    <= sub_wire5(52);
	sub_wire2(12, 53)    <= sub_wire5(53);
	sub_wire2(12, 54)    <= sub_wire5(54);
	sub_wire2(12, 55)    <= sub_wire5(55);
	sub_wire2(12, 56)    <= sub_wire5(56);
	sub_wire2(12, 57)    <= sub_wire5(57);
	sub_wire2(12, 58)    <= sub_wire5(58);
	sub_wire2(12, 59)    <= sub_wire5(59);
	sub_wire2(12, 60)    <= sub_wire5(60);
	sub_wire2(12, 61)    <= sub_wire5(61);
	sub_wire2(12, 62)    <= sub_wire5(62);
	sub_wire2(12, 63)    <= sub_wire5(63);
	sub_wire2(12, 64)    <= sub_wire5(64);
	sub_wire2(12, 65)    <= sub_wire5(65);
	sub_wire2(12, 66)    <= sub_wire5(66);
	sub_wire2(12, 67)    <= sub_wire5(67);
	sub_wire2(12, 68)    <= sub_wire5(68);
	sub_wire2(12, 69)    <= sub_wire5(69);
	sub_wire2(12, 70)    <= sub_wire5(70);
	sub_wire2(12, 71)    <= sub_wire5(71);
	sub_wire2(12, 72)    <= sub_wire5(72);
	sub_wire2(12, 73)    <= sub_wire5(73);
	sub_wire2(12, 74)    <= sub_wire5(74);
	sub_wire2(12, 75)    <= sub_wire5(75);
	sub_wire2(12, 76)    <= sub_wire5(76);
	sub_wire2(12, 77)    <= sub_wire5(77);
	sub_wire2(12, 78)    <= sub_wire5(78);
	sub_wire2(12, 79)    <= sub_wire5(79);
	sub_wire2(12, 80)    <= sub_wire5(80);
	sub_wire2(12, 81)    <= sub_wire5(81);
	sub_wire2(12, 82)    <= sub_wire5(82);
	sub_wire2(12, 83)    <= sub_wire5(83);
	sub_wire2(12, 84)    <= sub_wire5(84);
	sub_wire2(12, 85)    <= sub_wire5(85);
	sub_wire2(12, 86)    <= sub_wire5(86);
	sub_wire2(12, 87)    <= sub_wire5(87);
	sub_wire2(12, 88)    <= sub_wire5(88);
	sub_wire2(12, 89)    <= sub_wire5(89);
	sub_wire2(12, 90)    <= sub_wire5(90);
	sub_wire2(12, 91)    <= sub_wire5(91);
	sub_wire2(12, 92)    <= sub_wire5(92);
	sub_wire2(12, 93)    <= sub_wire5(93);
	sub_wire2(12, 94)    <= sub_wire5(94);
	sub_wire2(12, 95)    <= sub_wire5(95);
	sub_wire2(12, 96)    <= sub_wire5(96);
	sub_wire2(12, 97)    <= sub_wire5(97);
	sub_wire2(12, 98)    <= sub_wire5(98);
	sub_wire2(12, 99)    <= sub_wire5(99);
	sub_wire2(12, 100)    <= sub_wire5(100);
	sub_wire2(12, 101)    <= sub_wire5(101);
	sub_wire2(12, 102)    <= sub_wire5(102);
	sub_wire2(12, 103)    <= sub_wire5(103);
	sub_wire2(12, 104)    <= sub_wire5(104);
	sub_wire2(12, 105)    <= sub_wire5(105);
	sub_wire2(12, 106)    <= sub_wire5(106);
	sub_wire2(12, 107)    <= sub_wire5(107);
	sub_wire2(12, 108)    <= sub_wire5(108);
	sub_wire2(12, 109)    <= sub_wire5(109);
	sub_wire2(12, 110)    <= sub_wire5(110);
	sub_wire2(12, 111)    <= sub_wire5(111);
	sub_wire2(12, 112)    <= sub_wire5(112);
	sub_wire2(12, 113)    <= sub_wire5(113);
	sub_wire2(12, 114)    <= sub_wire5(114);
	sub_wire2(12, 115)    <= sub_wire5(115);
	sub_wire2(12, 116)    <= sub_wire5(116);
	sub_wire2(12, 117)    <= sub_wire5(117);
	sub_wire2(12, 118)    <= sub_wire5(118);
	sub_wire2(12, 119)    <= sub_wire5(119);
	sub_wire2(12, 120)    <= sub_wire5(120);
	sub_wire2(12, 121)    <= sub_wire5(121);
	sub_wire2(12, 122)    <= sub_wire5(122);
	sub_wire2(12, 123)    <= sub_wire5(123);
	sub_wire2(12, 124)    <= sub_wire5(124);
	sub_wire2(12, 125)    <= sub_wire5(125);
	sub_wire2(12, 126)    <= sub_wire5(126);
	sub_wire2(12, 127)    <= sub_wire5(127);
	sub_wire2(11, 0)    <= sub_wire6(0);
	sub_wire2(11, 1)    <= sub_wire6(1);
	sub_wire2(11, 2)    <= sub_wire6(2);
	sub_wire2(11, 3)    <= sub_wire6(3);
	sub_wire2(11, 4)    <= sub_wire6(4);
	sub_wire2(11, 5)    <= sub_wire6(5);
	sub_wire2(11, 6)    <= sub_wire6(6);
	sub_wire2(11, 7)    <= sub_wire6(7);
	sub_wire2(11, 8)    <= sub_wire6(8);
	sub_wire2(11, 9)    <= sub_wire6(9);
	sub_wire2(11, 10)    <= sub_wire6(10);
	sub_wire2(11, 11)    <= sub_wire6(11);
	sub_wire2(11, 12)    <= sub_wire6(12);
	sub_wire2(11, 13)    <= sub_wire6(13);
	sub_wire2(11, 14)    <= sub_wire6(14);
	sub_wire2(11, 15)    <= sub_wire6(15);
	sub_wire2(11, 16)    <= sub_wire6(16);
	sub_wire2(11, 17)    <= sub_wire6(17);
	sub_wire2(11, 18)    <= sub_wire6(18);
	sub_wire2(11, 19)    <= sub_wire6(19);
	sub_wire2(11, 20)    <= sub_wire6(20);
	sub_wire2(11, 21)    <= sub_wire6(21);
	sub_wire2(11, 22)    <= sub_wire6(22);
	sub_wire2(11, 23)    <= sub_wire6(23);
	sub_wire2(11, 24)    <= sub_wire6(24);
	sub_wire2(11, 25)    <= sub_wire6(25);
	sub_wire2(11, 26)    <= sub_wire6(26);
	sub_wire2(11, 27)    <= sub_wire6(27);
	sub_wire2(11, 28)    <= sub_wire6(28);
	sub_wire2(11, 29)    <= sub_wire6(29);
	sub_wire2(11, 30)    <= sub_wire6(30);
	sub_wire2(11, 31)    <= sub_wire6(31);
	sub_wire2(11, 32)    <= sub_wire6(32);
	sub_wire2(11, 33)    <= sub_wire6(33);
	sub_wire2(11, 34)    <= sub_wire6(34);
	sub_wire2(11, 35)    <= sub_wire6(35);
	sub_wire2(11, 36)    <= sub_wire6(36);
	sub_wire2(11, 37)    <= sub_wire6(37);
	sub_wire2(11, 38)    <= sub_wire6(38);
	sub_wire2(11, 39)    <= sub_wire6(39);
	sub_wire2(11, 40)    <= sub_wire6(40);
	sub_wire2(11, 41)    <= sub_wire6(41);
	sub_wire2(11, 42)    <= sub_wire6(42);
	sub_wire2(11, 43)    <= sub_wire6(43);
	sub_wire2(11, 44)    <= sub_wire6(44);
	sub_wire2(11, 45)    <= sub_wire6(45);
	sub_wire2(11, 46)    <= sub_wire6(46);
	sub_wire2(11, 47)    <= sub_wire6(47);
	sub_wire2(11, 48)    <= sub_wire6(48);
	sub_wire2(11, 49)    <= sub_wire6(49);
	sub_wire2(11, 50)    <= sub_wire6(50);
	sub_wire2(11, 51)    <= sub_wire6(51);
	sub_wire2(11, 52)    <= sub_wire6(52);
	sub_wire2(11, 53)    <= sub_wire6(53);
	sub_wire2(11, 54)    <= sub_wire6(54);
	sub_wire2(11, 55)    <= sub_wire6(55);
	sub_wire2(11, 56)    <= sub_wire6(56);
	sub_wire2(11, 57)    <= sub_wire6(57);
	sub_wire2(11, 58)    <= sub_wire6(58);
	sub_wire2(11, 59)    <= sub_wire6(59);
	sub_wire2(11, 60)    <= sub_wire6(60);
	sub_wire2(11, 61)    <= sub_wire6(61);
	sub_wire2(11, 62)    <= sub_wire6(62);
	sub_wire2(11, 63)    <= sub_wire6(63);
	sub_wire2(11, 64)    <= sub_wire6(64);
	sub_wire2(11, 65)    <= sub_wire6(65);
	sub_wire2(11, 66)    <= sub_wire6(66);
	sub_wire2(11, 67)    <= sub_wire6(67);
	sub_wire2(11, 68)    <= sub_wire6(68);
	sub_wire2(11, 69)    <= sub_wire6(69);
	sub_wire2(11, 70)    <= sub_wire6(70);
	sub_wire2(11, 71)    <= sub_wire6(71);
	sub_wire2(11, 72)    <= sub_wire6(72);
	sub_wire2(11, 73)    <= sub_wire6(73);
	sub_wire2(11, 74)    <= sub_wire6(74);
	sub_wire2(11, 75)    <= sub_wire6(75);
	sub_wire2(11, 76)    <= sub_wire6(76);
	sub_wire2(11, 77)    <= sub_wire6(77);
	sub_wire2(11, 78)    <= sub_wire6(78);
	sub_wire2(11, 79)    <= sub_wire6(79);
	sub_wire2(11, 80)    <= sub_wire6(80);
	sub_wire2(11, 81)    <= sub_wire6(81);
	sub_wire2(11, 82)    <= sub_wire6(82);
	sub_wire2(11, 83)    <= sub_wire6(83);
	sub_wire2(11, 84)    <= sub_wire6(84);
	sub_wire2(11, 85)    <= sub_wire6(85);
	sub_wire2(11, 86)    <= sub_wire6(86);
	sub_wire2(11, 87)    <= sub_wire6(87);
	sub_wire2(11, 88)    <= sub_wire6(88);
	sub_wire2(11, 89)    <= sub_wire6(89);
	sub_wire2(11, 90)    <= sub_wire6(90);
	sub_wire2(11, 91)    <= sub_wire6(91);
	sub_wire2(11, 92)    <= sub_wire6(92);
	sub_wire2(11, 93)    <= sub_wire6(93);
	sub_wire2(11, 94)    <= sub_wire6(94);
	sub_wire2(11, 95)    <= sub_wire6(95);
	sub_wire2(11, 96)    <= sub_wire6(96);
	sub_wire2(11, 97)    <= sub_wire6(97);
	sub_wire2(11, 98)    <= sub_wire6(98);
	sub_wire2(11, 99)    <= sub_wire6(99);
	sub_wire2(11, 100)    <= sub_wire6(100);
	sub_wire2(11, 101)    <= sub_wire6(101);
	sub_wire2(11, 102)    <= sub_wire6(102);
	sub_wire2(11, 103)    <= sub_wire6(103);
	sub_wire2(11, 104)    <= sub_wire6(104);
	sub_wire2(11, 105)    <= sub_wire6(105);
	sub_wire2(11, 106)    <= sub_wire6(106);
	sub_wire2(11, 107)    <= sub_wire6(107);
	sub_wire2(11, 108)    <= sub_wire6(108);
	sub_wire2(11, 109)    <= sub_wire6(109);
	sub_wire2(11, 110)    <= sub_wire6(110);
	sub_wire2(11, 111)    <= sub_wire6(111);
	sub_wire2(11, 112)    <= sub_wire6(112);
	sub_wire2(11, 113)    <= sub_wire6(113);
	sub_wire2(11, 114)    <= sub_wire6(114);
	sub_wire2(11, 115)    <= sub_wire6(115);
	sub_wire2(11, 116)    <= sub_wire6(116);
	sub_wire2(11, 117)    <= sub_wire6(117);
	sub_wire2(11, 118)    <= sub_wire6(118);
	sub_wire2(11, 119)    <= sub_wire6(119);
	sub_wire2(11, 120)    <= sub_wire6(120);
	sub_wire2(11, 121)    <= sub_wire6(121);
	sub_wire2(11, 122)    <= sub_wire6(122);
	sub_wire2(11, 123)    <= sub_wire6(123);
	sub_wire2(11, 124)    <= sub_wire6(124);
	sub_wire2(11, 125)    <= sub_wire6(125);
	sub_wire2(11, 126)    <= sub_wire6(126);
	sub_wire2(11, 127)    <= sub_wire6(127);
	sub_wire2(10, 0)    <= sub_wire7(0);
	sub_wire2(10, 1)    <= sub_wire7(1);
	sub_wire2(10, 2)    <= sub_wire7(2);
	sub_wire2(10, 3)    <= sub_wire7(3);
	sub_wire2(10, 4)    <= sub_wire7(4);
	sub_wire2(10, 5)    <= sub_wire7(5);
	sub_wire2(10, 6)    <= sub_wire7(6);
	sub_wire2(10, 7)    <= sub_wire7(7);
	sub_wire2(10, 8)    <= sub_wire7(8);
	sub_wire2(10, 9)    <= sub_wire7(9);
	sub_wire2(10, 10)    <= sub_wire7(10);
	sub_wire2(10, 11)    <= sub_wire7(11);
	sub_wire2(10, 12)    <= sub_wire7(12);
	sub_wire2(10, 13)    <= sub_wire7(13);
	sub_wire2(10, 14)    <= sub_wire7(14);
	sub_wire2(10, 15)    <= sub_wire7(15);
	sub_wire2(10, 16)    <= sub_wire7(16);
	sub_wire2(10, 17)    <= sub_wire7(17);
	sub_wire2(10, 18)    <= sub_wire7(18);
	sub_wire2(10, 19)    <= sub_wire7(19);
	sub_wire2(10, 20)    <= sub_wire7(20);
	sub_wire2(10, 21)    <= sub_wire7(21);
	sub_wire2(10, 22)    <= sub_wire7(22);
	sub_wire2(10, 23)    <= sub_wire7(23);
	sub_wire2(10, 24)    <= sub_wire7(24);
	sub_wire2(10, 25)    <= sub_wire7(25);
	sub_wire2(10, 26)    <= sub_wire7(26);
	sub_wire2(10, 27)    <= sub_wire7(27);
	sub_wire2(10, 28)    <= sub_wire7(28);
	sub_wire2(10, 29)    <= sub_wire7(29);
	sub_wire2(10, 30)    <= sub_wire7(30);
	sub_wire2(10, 31)    <= sub_wire7(31);
	sub_wire2(10, 32)    <= sub_wire7(32);
	sub_wire2(10, 33)    <= sub_wire7(33);
	sub_wire2(10, 34)    <= sub_wire7(34);
	sub_wire2(10, 35)    <= sub_wire7(35);
	sub_wire2(10, 36)    <= sub_wire7(36);
	sub_wire2(10, 37)    <= sub_wire7(37);
	sub_wire2(10, 38)    <= sub_wire7(38);
	sub_wire2(10, 39)    <= sub_wire7(39);
	sub_wire2(10, 40)    <= sub_wire7(40);
	sub_wire2(10, 41)    <= sub_wire7(41);
	sub_wire2(10, 42)    <= sub_wire7(42);
	sub_wire2(10, 43)    <= sub_wire7(43);
	sub_wire2(10, 44)    <= sub_wire7(44);
	sub_wire2(10, 45)    <= sub_wire7(45);
	sub_wire2(10, 46)    <= sub_wire7(46);
	sub_wire2(10, 47)    <= sub_wire7(47);
	sub_wire2(10, 48)    <= sub_wire7(48);
	sub_wire2(10, 49)    <= sub_wire7(49);
	sub_wire2(10, 50)    <= sub_wire7(50);
	sub_wire2(10, 51)    <= sub_wire7(51);
	sub_wire2(10, 52)    <= sub_wire7(52);
	sub_wire2(10, 53)    <= sub_wire7(53);
	sub_wire2(10, 54)    <= sub_wire7(54);
	sub_wire2(10, 55)    <= sub_wire7(55);
	sub_wire2(10, 56)    <= sub_wire7(56);
	sub_wire2(10, 57)    <= sub_wire7(57);
	sub_wire2(10, 58)    <= sub_wire7(58);
	sub_wire2(10, 59)    <= sub_wire7(59);
	sub_wire2(10, 60)    <= sub_wire7(60);
	sub_wire2(10, 61)    <= sub_wire7(61);
	sub_wire2(10, 62)    <= sub_wire7(62);
	sub_wire2(10, 63)    <= sub_wire7(63);
	sub_wire2(10, 64)    <= sub_wire7(64);
	sub_wire2(10, 65)    <= sub_wire7(65);
	sub_wire2(10, 66)    <= sub_wire7(66);
	sub_wire2(10, 67)    <= sub_wire7(67);
	sub_wire2(10, 68)    <= sub_wire7(68);
	sub_wire2(10, 69)    <= sub_wire7(69);
	sub_wire2(10, 70)    <= sub_wire7(70);
	sub_wire2(10, 71)    <= sub_wire7(71);
	sub_wire2(10, 72)    <= sub_wire7(72);
	sub_wire2(10, 73)    <= sub_wire7(73);
	sub_wire2(10, 74)    <= sub_wire7(74);
	sub_wire2(10, 75)    <= sub_wire7(75);
	sub_wire2(10, 76)    <= sub_wire7(76);
	sub_wire2(10, 77)    <= sub_wire7(77);
	sub_wire2(10, 78)    <= sub_wire7(78);
	sub_wire2(10, 79)    <= sub_wire7(79);
	sub_wire2(10, 80)    <= sub_wire7(80);
	sub_wire2(10, 81)    <= sub_wire7(81);
	sub_wire2(10, 82)    <= sub_wire7(82);
	sub_wire2(10, 83)    <= sub_wire7(83);
	sub_wire2(10, 84)    <= sub_wire7(84);
	sub_wire2(10, 85)    <= sub_wire7(85);
	sub_wire2(10, 86)    <= sub_wire7(86);
	sub_wire2(10, 87)    <= sub_wire7(87);
	sub_wire2(10, 88)    <= sub_wire7(88);
	sub_wire2(10, 89)    <= sub_wire7(89);
	sub_wire2(10, 90)    <= sub_wire7(90);
	sub_wire2(10, 91)    <= sub_wire7(91);
	sub_wire2(10, 92)    <= sub_wire7(92);
	sub_wire2(10, 93)    <= sub_wire7(93);
	sub_wire2(10, 94)    <= sub_wire7(94);
	sub_wire2(10, 95)    <= sub_wire7(95);
	sub_wire2(10, 96)    <= sub_wire7(96);
	sub_wire2(10, 97)    <= sub_wire7(97);
	sub_wire2(10, 98)    <= sub_wire7(98);
	sub_wire2(10, 99)    <= sub_wire7(99);
	sub_wire2(10, 100)    <= sub_wire7(100);
	sub_wire2(10, 101)    <= sub_wire7(101);
	sub_wire2(10, 102)    <= sub_wire7(102);
	sub_wire2(10, 103)    <= sub_wire7(103);
	sub_wire2(10, 104)    <= sub_wire7(104);
	sub_wire2(10, 105)    <= sub_wire7(105);
	sub_wire2(10, 106)    <= sub_wire7(106);
	sub_wire2(10, 107)    <= sub_wire7(107);
	sub_wire2(10, 108)    <= sub_wire7(108);
	sub_wire2(10, 109)    <= sub_wire7(109);
	sub_wire2(10, 110)    <= sub_wire7(110);
	sub_wire2(10, 111)    <= sub_wire7(111);
	sub_wire2(10, 112)    <= sub_wire7(112);
	sub_wire2(10, 113)    <= sub_wire7(113);
	sub_wire2(10, 114)    <= sub_wire7(114);
	sub_wire2(10, 115)    <= sub_wire7(115);
	sub_wire2(10, 116)    <= sub_wire7(116);
	sub_wire2(10, 117)    <= sub_wire7(117);
	sub_wire2(10, 118)    <= sub_wire7(118);
	sub_wire2(10, 119)    <= sub_wire7(119);
	sub_wire2(10, 120)    <= sub_wire7(120);
	sub_wire2(10, 121)    <= sub_wire7(121);
	sub_wire2(10, 122)    <= sub_wire7(122);
	sub_wire2(10, 123)    <= sub_wire7(123);
	sub_wire2(10, 124)    <= sub_wire7(124);
	sub_wire2(10, 125)    <= sub_wire7(125);
	sub_wire2(10, 126)    <= sub_wire7(126);
	sub_wire2(10, 127)    <= sub_wire7(127);
	sub_wire2(9, 0)    <= sub_wire8(0);
	sub_wire2(9, 1)    <= sub_wire8(1);
	sub_wire2(9, 2)    <= sub_wire8(2);
	sub_wire2(9, 3)    <= sub_wire8(3);
	sub_wire2(9, 4)    <= sub_wire8(4);
	sub_wire2(9, 5)    <= sub_wire8(5);
	sub_wire2(9, 6)    <= sub_wire8(6);
	sub_wire2(9, 7)    <= sub_wire8(7);
	sub_wire2(9, 8)    <= sub_wire8(8);
	sub_wire2(9, 9)    <= sub_wire8(9);
	sub_wire2(9, 10)    <= sub_wire8(10);
	sub_wire2(9, 11)    <= sub_wire8(11);
	sub_wire2(9, 12)    <= sub_wire8(12);
	sub_wire2(9, 13)    <= sub_wire8(13);
	sub_wire2(9, 14)    <= sub_wire8(14);
	sub_wire2(9, 15)    <= sub_wire8(15);
	sub_wire2(9, 16)    <= sub_wire8(16);
	sub_wire2(9, 17)    <= sub_wire8(17);
	sub_wire2(9, 18)    <= sub_wire8(18);
	sub_wire2(9, 19)    <= sub_wire8(19);
	sub_wire2(9, 20)    <= sub_wire8(20);
	sub_wire2(9, 21)    <= sub_wire8(21);
	sub_wire2(9, 22)    <= sub_wire8(22);
	sub_wire2(9, 23)    <= sub_wire8(23);
	sub_wire2(9, 24)    <= sub_wire8(24);
	sub_wire2(9, 25)    <= sub_wire8(25);
	sub_wire2(9, 26)    <= sub_wire8(26);
	sub_wire2(9, 27)    <= sub_wire8(27);
	sub_wire2(9, 28)    <= sub_wire8(28);
	sub_wire2(9, 29)    <= sub_wire8(29);
	sub_wire2(9, 30)    <= sub_wire8(30);
	sub_wire2(9, 31)    <= sub_wire8(31);
	sub_wire2(9, 32)    <= sub_wire8(32);
	sub_wire2(9, 33)    <= sub_wire8(33);
	sub_wire2(9, 34)    <= sub_wire8(34);
	sub_wire2(9, 35)    <= sub_wire8(35);
	sub_wire2(9, 36)    <= sub_wire8(36);
	sub_wire2(9, 37)    <= sub_wire8(37);
	sub_wire2(9, 38)    <= sub_wire8(38);
	sub_wire2(9, 39)    <= sub_wire8(39);
	sub_wire2(9, 40)    <= sub_wire8(40);
	sub_wire2(9, 41)    <= sub_wire8(41);
	sub_wire2(9, 42)    <= sub_wire8(42);
	sub_wire2(9, 43)    <= sub_wire8(43);
	sub_wire2(9, 44)    <= sub_wire8(44);
	sub_wire2(9, 45)    <= sub_wire8(45);
	sub_wire2(9, 46)    <= sub_wire8(46);
	sub_wire2(9, 47)    <= sub_wire8(47);
	sub_wire2(9, 48)    <= sub_wire8(48);
	sub_wire2(9, 49)    <= sub_wire8(49);
	sub_wire2(9, 50)    <= sub_wire8(50);
	sub_wire2(9, 51)    <= sub_wire8(51);
	sub_wire2(9, 52)    <= sub_wire8(52);
	sub_wire2(9, 53)    <= sub_wire8(53);
	sub_wire2(9, 54)    <= sub_wire8(54);
	sub_wire2(9, 55)    <= sub_wire8(55);
	sub_wire2(9, 56)    <= sub_wire8(56);
	sub_wire2(9, 57)    <= sub_wire8(57);
	sub_wire2(9, 58)    <= sub_wire8(58);
	sub_wire2(9, 59)    <= sub_wire8(59);
	sub_wire2(9, 60)    <= sub_wire8(60);
	sub_wire2(9, 61)    <= sub_wire8(61);
	sub_wire2(9, 62)    <= sub_wire8(62);
	sub_wire2(9, 63)    <= sub_wire8(63);
	sub_wire2(9, 64)    <= sub_wire8(64);
	sub_wire2(9, 65)    <= sub_wire8(65);
	sub_wire2(9, 66)    <= sub_wire8(66);
	sub_wire2(9, 67)    <= sub_wire8(67);
	sub_wire2(9, 68)    <= sub_wire8(68);
	sub_wire2(9, 69)    <= sub_wire8(69);
	sub_wire2(9, 70)    <= sub_wire8(70);
	sub_wire2(9, 71)    <= sub_wire8(71);
	sub_wire2(9, 72)    <= sub_wire8(72);
	sub_wire2(9, 73)    <= sub_wire8(73);
	sub_wire2(9, 74)    <= sub_wire8(74);
	sub_wire2(9, 75)    <= sub_wire8(75);
	sub_wire2(9, 76)    <= sub_wire8(76);
	sub_wire2(9, 77)    <= sub_wire8(77);
	sub_wire2(9, 78)    <= sub_wire8(78);
	sub_wire2(9, 79)    <= sub_wire8(79);
	sub_wire2(9, 80)    <= sub_wire8(80);
	sub_wire2(9, 81)    <= sub_wire8(81);
	sub_wire2(9, 82)    <= sub_wire8(82);
	sub_wire2(9, 83)    <= sub_wire8(83);
	sub_wire2(9, 84)    <= sub_wire8(84);
	sub_wire2(9, 85)    <= sub_wire8(85);
	sub_wire2(9, 86)    <= sub_wire8(86);
	sub_wire2(9, 87)    <= sub_wire8(87);
	sub_wire2(9, 88)    <= sub_wire8(88);
	sub_wire2(9, 89)    <= sub_wire8(89);
	sub_wire2(9, 90)    <= sub_wire8(90);
	sub_wire2(9, 91)    <= sub_wire8(91);
	sub_wire2(9, 92)    <= sub_wire8(92);
	sub_wire2(9, 93)    <= sub_wire8(93);
	sub_wire2(9, 94)    <= sub_wire8(94);
	sub_wire2(9, 95)    <= sub_wire8(95);
	sub_wire2(9, 96)    <= sub_wire8(96);
	sub_wire2(9, 97)    <= sub_wire8(97);
	sub_wire2(9, 98)    <= sub_wire8(98);
	sub_wire2(9, 99)    <= sub_wire8(99);
	sub_wire2(9, 100)    <= sub_wire8(100);
	sub_wire2(9, 101)    <= sub_wire8(101);
	sub_wire2(9, 102)    <= sub_wire8(102);
	sub_wire2(9, 103)    <= sub_wire8(103);
	sub_wire2(9, 104)    <= sub_wire8(104);
	sub_wire2(9, 105)    <= sub_wire8(105);
	sub_wire2(9, 106)    <= sub_wire8(106);
	sub_wire2(9, 107)    <= sub_wire8(107);
	sub_wire2(9, 108)    <= sub_wire8(108);
	sub_wire2(9, 109)    <= sub_wire8(109);
	sub_wire2(9, 110)    <= sub_wire8(110);
	sub_wire2(9, 111)    <= sub_wire8(111);
	sub_wire2(9, 112)    <= sub_wire8(112);
	sub_wire2(9, 113)    <= sub_wire8(113);
	sub_wire2(9, 114)    <= sub_wire8(114);
	sub_wire2(9, 115)    <= sub_wire8(115);
	sub_wire2(9, 116)    <= sub_wire8(116);
	sub_wire2(9, 117)    <= sub_wire8(117);
	sub_wire2(9, 118)    <= sub_wire8(118);
	sub_wire2(9, 119)    <= sub_wire8(119);
	sub_wire2(9, 120)    <= sub_wire8(120);
	sub_wire2(9, 121)    <= sub_wire8(121);
	sub_wire2(9, 122)    <= sub_wire8(122);
	sub_wire2(9, 123)    <= sub_wire8(123);
	sub_wire2(9, 124)    <= sub_wire8(124);
	sub_wire2(9, 125)    <= sub_wire8(125);
	sub_wire2(9, 126)    <= sub_wire8(126);
	sub_wire2(9, 127)    <= sub_wire8(127);
	sub_wire2(8, 0)    <= sub_wire9(0);
	sub_wire2(8, 1)    <= sub_wire9(1);
	sub_wire2(8, 2)    <= sub_wire9(2);
	sub_wire2(8, 3)    <= sub_wire9(3);
	sub_wire2(8, 4)    <= sub_wire9(4);
	sub_wire2(8, 5)    <= sub_wire9(5);
	sub_wire2(8, 6)    <= sub_wire9(6);
	sub_wire2(8, 7)    <= sub_wire9(7);
	sub_wire2(8, 8)    <= sub_wire9(8);
	sub_wire2(8, 9)    <= sub_wire9(9);
	sub_wire2(8, 10)    <= sub_wire9(10);
	sub_wire2(8, 11)    <= sub_wire9(11);
	sub_wire2(8, 12)    <= sub_wire9(12);
	sub_wire2(8, 13)    <= sub_wire9(13);
	sub_wire2(8, 14)    <= sub_wire9(14);
	sub_wire2(8, 15)    <= sub_wire9(15);
	sub_wire2(8, 16)    <= sub_wire9(16);
	sub_wire2(8, 17)    <= sub_wire9(17);
	sub_wire2(8, 18)    <= sub_wire9(18);
	sub_wire2(8, 19)    <= sub_wire9(19);
	sub_wire2(8, 20)    <= sub_wire9(20);
	sub_wire2(8, 21)    <= sub_wire9(21);
	sub_wire2(8, 22)    <= sub_wire9(22);
	sub_wire2(8, 23)    <= sub_wire9(23);
	sub_wire2(8, 24)    <= sub_wire9(24);
	sub_wire2(8, 25)    <= sub_wire9(25);
	sub_wire2(8, 26)    <= sub_wire9(26);
	sub_wire2(8, 27)    <= sub_wire9(27);
	sub_wire2(8, 28)    <= sub_wire9(28);
	sub_wire2(8, 29)    <= sub_wire9(29);
	sub_wire2(8, 30)    <= sub_wire9(30);
	sub_wire2(8, 31)    <= sub_wire9(31);
	sub_wire2(8, 32)    <= sub_wire9(32);
	sub_wire2(8, 33)    <= sub_wire9(33);
	sub_wire2(8, 34)    <= sub_wire9(34);
	sub_wire2(8, 35)    <= sub_wire9(35);
	sub_wire2(8, 36)    <= sub_wire9(36);
	sub_wire2(8, 37)    <= sub_wire9(37);
	sub_wire2(8, 38)    <= sub_wire9(38);
	sub_wire2(8, 39)    <= sub_wire9(39);
	sub_wire2(8, 40)    <= sub_wire9(40);
	sub_wire2(8, 41)    <= sub_wire9(41);
	sub_wire2(8, 42)    <= sub_wire9(42);
	sub_wire2(8, 43)    <= sub_wire9(43);
	sub_wire2(8, 44)    <= sub_wire9(44);
	sub_wire2(8, 45)    <= sub_wire9(45);
	sub_wire2(8, 46)    <= sub_wire9(46);
	sub_wire2(8, 47)    <= sub_wire9(47);
	sub_wire2(8, 48)    <= sub_wire9(48);
	sub_wire2(8, 49)    <= sub_wire9(49);
	sub_wire2(8, 50)    <= sub_wire9(50);
	sub_wire2(8, 51)    <= sub_wire9(51);
	sub_wire2(8, 52)    <= sub_wire9(52);
	sub_wire2(8, 53)    <= sub_wire9(53);
	sub_wire2(8, 54)    <= sub_wire9(54);
	sub_wire2(8, 55)    <= sub_wire9(55);
	sub_wire2(8, 56)    <= sub_wire9(56);
	sub_wire2(8, 57)    <= sub_wire9(57);
	sub_wire2(8, 58)    <= sub_wire9(58);
	sub_wire2(8, 59)    <= sub_wire9(59);
	sub_wire2(8, 60)    <= sub_wire9(60);
	sub_wire2(8, 61)    <= sub_wire9(61);
	sub_wire2(8, 62)    <= sub_wire9(62);
	sub_wire2(8, 63)    <= sub_wire9(63);
	sub_wire2(8, 64)    <= sub_wire9(64);
	sub_wire2(8, 65)    <= sub_wire9(65);
	sub_wire2(8, 66)    <= sub_wire9(66);
	sub_wire2(8, 67)    <= sub_wire9(67);
	sub_wire2(8, 68)    <= sub_wire9(68);
	sub_wire2(8, 69)    <= sub_wire9(69);
	sub_wire2(8, 70)    <= sub_wire9(70);
	sub_wire2(8, 71)    <= sub_wire9(71);
	sub_wire2(8, 72)    <= sub_wire9(72);
	sub_wire2(8, 73)    <= sub_wire9(73);
	sub_wire2(8, 74)    <= sub_wire9(74);
	sub_wire2(8, 75)    <= sub_wire9(75);
	sub_wire2(8, 76)    <= sub_wire9(76);
	sub_wire2(8, 77)    <= sub_wire9(77);
	sub_wire2(8, 78)    <= sub_wire9(78);
	sub_wire2(8, 79)    <= sub_wire9(79);
	sub_wire2(8, 80)    <= sub_wire9(80);
	sub_wire2(8, 81)    <= sub_wire9(81);
	sub_wire2(8, 82)    <= sub_wire9(82);
	sub_wire2(8, 83)    <= sub_wire9(83);
	sub_wire2(8, 84)    <= sub_wire9(84);
	sub_wire2(8, 85)    <= sub_wire9(85);
	sub_wire2(8, 86)    <= sub_wire9(86);
	sub_wire2(8, 87)    <= sub_wire9(87);
	sub_wire2(8, 88)    <= sub_wire9(88);
	sub_wire2(8, 89)    <= sub_wire9(89);
	sub_wire2(8, 90)    <= sub_wire9(90);
	sub_wire2(8, 91)    <= sub_wire9(91);
	sub_wire2(8, 92)    <= sub_wire9(92);
	sub_wire2(8, 93)    <= sub_wire9(93);
	sub_wire2(8, 94)    <= sub_wire9(94);
	sub_wire2(8, 95)    <= sub_wire9(95);
	sub_wire2(8, 96)    <= sub_wire9(96);
	sub_wire2(8, 97)    <= sub_wire9(97);
	sub_wire2(8, 98)    <= sub_wire9(98);
	sub_wire2(8, 99)    <= sub_wire9(99);
	sub_wire2(8, 100)    <= sub_wire9(100);
	sub_wire2(8, 101)    <= sub_wire9(101);
	sub_wire2(8, 102)    <= sub_wire9(102);
	sub_wire2(8, 103)    <= sub_wire9(103);
	sub_wire2(8, 104)    <= sub_wire9(104);
	sub_wire2(8, 105)    <= sub_wire9(105);
	sub_wire2(8, 106)    <= sub_wire9(106);
	sub_wire2(8, 107)    <= sub_wire9(107);
	sub_wire2(8, 108)    <= sub_wire9(108);
	sub_wire2(8, 109)    <= sub_wire9(109);
	sub_wire2(8, 110)    <= sub_wire9(110);
	sub_wire2(8, 111)    <= sub_wire9(111);
	sub_wire2(8, 112)    <= sub_wire9(112);
	sub_wire2(8, 113)    <= sub_wire9(113);
	sub_wire2(8, 114)    <= sub_wire9(114);
	sub_wire2(8, 115)    <= sub_wire9(115);
	sub_wire2(8, 116)    <= sub_wire9(116);
	sub_wire2(8, 117)    <= sub_wire9(117);
	sub_wire2(8, 118)    <= sub_wire9(118);
	sub_wire2(8, 119)    <= sub_wire9(119);
	sub_wire2(8, 120)    <= sub_wire9(120);
	sub_wire2(8, 121)    <= sub_wire9(121);
	sub_wire2(8, 122)    <= sub_wire9(122);
	sub_wire2(8, 123)    <= sub_wire9(123);
	sub_wire2(8, 124)    <= sub_wire9(124);
	sub_wire2(8, 125)    <= sub_wire9(125);
	sub_wire2(8, 126)    <= sub_wire9(126);
	sub_wire2(8, 127)    <= sub_wire9(127);
	sub_wire2(7, 0)    <= sub_wire10(0);
	sub_wire2(7, 1)    <= sub_wire10(1);
	sub_wire2(7, 2)    <= sub_wire10(2);
	sub_wire2(7, 3)    <= sub_wire10(3);
	sub_wire2(7, 4)    <= sub_wire10(4);
	sub_wire2(7, 5)    <= sub_wire10(5);
	sub_wire2(7, 6)    <= sub_wire10(6);
	sub_wire2(7, 7)    <= sub_wire10(7);
	sub_wire2(7, 8)    <= sub_wire10(8);
	sub_wire2(7, 9)    <= sub_wire10(9);
	sub_wire2(7, 10)    <= sub_wire10(10);
	sub_wire2(7, 11)    <= sub_wire10(11);
	sub_wire2(7, 12)    <= sub_wire10(12);
	sub_wire2(7, 13)    <= sub_wire10(13);
	sub_wire2(7, 14)    <= sub_wire10(14);
	sub_wire2(7, 15)    <= sub_wire10(15);
	sub_wire2(7, 16)    <= sub_wire10(16);
	sub_wire2(7, 17)    <= sub_wire10(17);
	sub_wire2(7, 18)    <= sub_wire10(18);
	sub_wire2(7, 19)    <= sub_wire10(19);
	sub_wire2(7, 20)    <= sub_wire10(20);
	sub_wire2(7, 21)    <= sub_wire10(21);
	sub_wire2(7, 22)    <= sub_wire10(22);
	sub_wire2(7, 23)    <= sub_wire10(23);
	sub_wire2(7, 24)    <= sub_wire10(24);
	sub_wire2(7, 25)    <= sub_wire10(25);
	sub_wire2(7, 26)    <= sub_wire10(26);
	sub_wire2(7, 27)    <= sub_wire10(27);
	sub_wire2(7, 28)    <= sub_wire10(28);
	sub_wire2(7, 29)    <= sub_wire10(29);
	sub_wire2(7, 30)    <= sub_wire10(30);
	sub_wire2(7, 31)    <= sub_wire10(31);
	sub_wire2(7, 32)    <= sub_wire10(32);
	sub_wire2(7, 33)    <= sub_wire10(33);
	sub_wire2(7, 34)    <= sub_wire10(34);
	sub_wire2(7, 35)    <= sub_wire10(35);
	sub_wire2(7, 36)    <= sub_wire10(36);
	sub_wire2(7, 37)    <= sub_wire10(37);
	sub_wire2(7, 38)    <= sub_wire10(38);
	sub_wire2(7, 39)    <= sub_wire10(39);
	sub_wire2(7, 40)    <= sub_wire10(40);
	sub_wire2(7, 41)    <= sub_wire10(41);
	sub_wire2(7, 42)    <= sub_wire10(42);
	sub_wire2(7, 43)    <= sub_wire10(43);
	sub_wire2(7, 44)    <= sub_wire10(44);
	sub_wire2(7, 45)    <= sub_wire10(45);
	sub_wire2(7, 46)    <= sub_wire10(46);
	sub_wire2(7, 47)    <= sub_wire10(47);
	sub_wire2(7, 48)    <= sub_wire10(48);
	sub_wire2(7, 49)    <= sub_wire10(49);
	sub_wire2(7, 50)    <= sub_wire10(50);
	sub_wire2(7, 51)    <= sub_wire10(51);
	sub_wire2(7, 52)    <= sub_wire10(52);
	sub_wire2(7, 53)    <= sub_wire10(53);
	sub_wire2(7, 54)    <= sub_wire10(54);
	sub_wire2(7, 55)    <= sub_wire10(55);
	sub_wire2(7, 56)    <= sub_wire10(56);
	sub_wire2(7, 57)    <= sub_wire10(57);
	sub_wire2(7, 58)    <= sub_wire10(58);
	sub_wire2(7, 59)    <= sub_wire10(59);
	sub_wire2(7, 60)    <= sub_wire10(60);
	sub_wire2(7, 61)    <= sub_wire10(61);
	sub_wire2(7, 62)    <= sub_wire10(62);
	sub_wire2(7, 63)    <= sub_wire10(63);
	sub_wire2(7, 64)    <= sub_wire10(64);
	sub_wire2(7, 65)    <= sub_wire10(65);
	sub_wire2(7, 66)    <= sub_wire10(66);
	sub_wire2(7, 67)    <= sub_wire10(67);
	sub_wire2(7, 68)    <= sub_wire10(68);
	sub_wire2(7, 69)    <= sub_wire10(69);
	sub_wire2(7, 70)    <= sub_wire10(70);
	sub_wire2(7, 71)    <= sub_wire10(71);
	sub_wire2(7, 72)    <= sub_wire10(72);
	sub_wire2(7, 73)    <= sub_wire10(73);
	sub_wire2(7, 74)    <= sub_wire10(74);
	sub_wire2(7, 75)    <= sub_wire10(75);
	sub_wire2(7, 76)    <= sub_wire10(76);
	sub_wire2(7, 77)    <= sub_wire10(77);
	sub_wire2(7, 78)    <= sub_wire10(78);
	sub_wire2(7, 79)    <= sub_wire10(79);
	sub_wire2(7, 80)    <= sub_wire10(80);
	sub_wire2(7, 81)    <= sub_wire10(81);
	sub_wire2(7, 82)    <= sub_wire10(82);
	sub_wire2(7, 83)    <= sub_wire10(83);
	sub_wire2(7, 84)    <= sub_wire10(84);
	sub_wire2(7, 85)    <= sub_wire10(85);
	sub_wire2(7, 86)    <= sub_wire10(86);
	sub_wire2(7, 87)    <= sub_wire10(87);
	sub_wire2(7, 88)    <= sub_wire10(88);
	sub_wire2(7, 89)    <= sub_wire10(89);
	sub_wire2(7, 90)    <= sub_wire10(90);
	sub_wire2(7, 91)    <= sub_wire10(91);
	sub_wire2(7, 92)    <= sub_wire10(92);
	sub_wire2(7, 93)    <= sub_wire10(93);
	sub_wire2(7, 94)    <= sub_wire10(94);
	sub_wire2(7, 95)    <= sub_wire10(95);
	sub_wire2(7, 96)    <= sub_wire10(96);
	sub_wire2(7, 97)    <= sub_wire10(97);
	sub_wire2(7, 98)    <= sub_wire10(98);
	sub_wire2(7, 99)    <= sub_wire10(99);
	sub_wire2(7, 100)    <= sub_wire10(100);
	sub_wire2(7, 101)    <= sub_wire10(101);
	sub_wire2(7, 102)    <= sub_wire10(102);
	sub_wire2(7, 103)    <= sub_wire10(103);
	sub_wire2(7, 104)    <= sub_wire10(104);
	sub_wire2(7, 105)    <= sub_wire10(105);
	sub_wire2(7, 106)    <= sub_wire10(106);
	sub_wire2(7, 107)    <= sub_wire10(107);
	sub_wire2(7, 108)    <= sub_wire10(108);
	sub_wire2(7, 109)    <= sub_wire10(109);
	sub_wire2(7, 110)    <= sub_wire10(110);
	sub_wire2(7, 111)    <= sub_wire10(111);
	sub_wire2(7, 112)    <= sub_wire10(112);
	sub_wire2(7, 113)    <= sub_wire10(113);
	sub_wire2(7, 114)    <= sub_wire10(114);
	sub_wire2(7, 115)    <= sub_wire10(115);
	sub_wire2(7, 116)    <= sub_wire10(116);
	sub_wire2(7, 117)    <= sub_wire10(117);
	sub_wire2(7, 118)    <= sub_wire10(118);
	sub_wire2(7, 119)    <= sub_wire10(119);
	sub_wire2(7, 120)    <= sub_wire10(120);
	sub_wire2(7, 121)    <= sub_wire10(121);
	sub_wire2(7, 122)    <= sub_wire10(122);
	sub_wire2(7, 123)    <= sub_wire10(123);
	sub_wire2(7, 124)    <= sub_wire10(124);
	sub_wire2(7, 125)    <= sub_wire10(125);
	sub_wire2(7, 126)    <= sub_wire10(126);
	sub_wire2(7, 127)    <= sub_wire10(127);
	sub_wire2(6, 0)    <= sub_wire11(0);
	sub_wire2(6, 1)    <= sub_wire11(1);
	sub_wire2(6, 2)    <= sub_wire11(2);
	sub_wire2(6, 3)    <= sub_wire11(3);
	sub_wire2(6, 4)    <= sub_wire11(4);
	sub_wire2(6, 5)    <= sub_wire11(5);
	sub_wire2(6, 6)    <= sub_wire11(6);
	sub_wire2(6, 7)    <= sub_wire11(7);
	sub_wire2(6, 8)    <= sub_wire11(8);
	sub_wire2(6, 9)    <= sub_wire11(9);
	sub_wire2(6, 10)    <= sub_wire11(10);
	sub_wire2(6, 11)    <= sub_wire11(11);
	sub_wire2(6, 12)    <= sub_wire11(12);
	sub_wire2(6, 13)    <= sub_wire11(13);
	sub_wire2(6, 14)    <= sub_wire11(14);
	sub_wire2(6, 15)    <= sub_wire11(15);
	sub_wire2(6, 16)    <= sub_wire11(16);
	sub_wire2(6, 17)    <= sub_wire11(17);
	sub_wire2(6, 18)    <= sub_wire11(18);
	sub_wire2(6, 19)    <= sub_wire11(19);
	sub_wire2(6, 20)    <= sub_wire11(20);
	sub_wire2(6, 21)    <= sub_wire11(21);
	sub_wire2(6, 22)    <= sub_wire11(22);
	sub_wire2(6, 23)    <= sub_wire11(23);
	sub_wire2(6, 24)    <= sub_wire11(24);
	sub_wire2(6, 25)    <= sub_wire11(25);
	sub_wire2(6, 26)    <= sub_wire11(26);
	sub_wire2(6, 27)    <= sub_wire11(27);
	sub_wire2(6, 28)    <= sub_wire11(28);
	sub_wire2(6, 29)    <= sub_wire11(29);
	sub_wire2(6, 30)    <= sub_wire11(30);
	sub_wire2(6, 31)    <= sub_wire11(31);
	sub_wire2(6, 32)    <= sub_wire11(32);
	sub_wire2(6, 33)    <= sub_wire11(33);
	sub_wire2(6, 34)    <= sub_wire11(34);
	sub_wire2(6, 35)    <= sub_wire11(35);
	sub_wire2(6, 36)    <= sub_wire11(36);
	sub_wire2(6, 37)    <= sub_wire11(37);
	sub_wire2(6, 38)    <= sub_wire11(38);
	sub_wire2(6, 39)    <= sub_wire11(39);
	sub_wire2(6, 40)    <= sub_wire11(40);
	sub_wire2(6, 41)    <= sub_wire11(41);
	sub_wire2(6, 42)    <= sub_wire11(42);
	sub_wire2(6, 43)    <= sub_wire11(43);
	sub_wire2(6, 44)    <= sub_wire11(44);
	sub_wire2(6, 45)    <= sub_wire11(45);
	sub_wire2(6, 46)    <= sub_wire11(46);
	sub_wire2(6, 47)    <= sub_wire11(47);
	sub_wire2(6, 48)    <= sub_wire11(48);
	sub_wire2(6, 49)    <= sub_wire11(49);
	sub_wire2(6, 50)    <= sub_wire11(50);
	sub_wire2(6, 51)    <= sub_wire11(51);
	sub_wire2(6, 52)    <= sub_wire11(52);
	sub_wire2(6, 53)    <= sub_wire11(53);
	sub_wire2(6, 54)    <= sub_wire11(54);
	sub_wire2(6, 55)    <= sub_wire11(55);
	sub_wire2(6, 56)    <= sub_wire11(56);
	sub_wire2(6, 57)    <= sub_wire11(57);
	sub_wire2(6, 58)    <= sub_wire11(58);
	sub_wire2(6, 59)    <= sub_wire11(59);
	sub_wire2(6, 60)    <= sub_wire11(60);
	sub_wire2(6, 61)    <= sub_wire11(61);
	sub_wire2(6, 62)    <= sub_wire11(62);
	sub_wire2(6, 63)    <= sub_wire11(63);
	sub_wire2(6, 64)    <= sub_wire11(64);
	sub_wire2(6, 65)    <= sub_wire11(65);
	sub_wire2(6, 66)    <= sub_wire11(66);
	sub_wire2(6, 67)    <= sub_wire11(67);
	sub_wire2(6, 68)    <= sub_wire11(68);
	sub_wire2(6, 69)    <= sub_wire11(69);
	sub_wire2(6, 70)    <= sub_wire11(70);
	sub_wire2(6, 71)    <= sub_wire11(71);
	sub_wire2(6, 72)    <= sub_wire11(72);
	sub_wire2(6, 73)    <= sub_wire11(73);
	sub_wire2(6, 74)    <= sub_wire11(74);
	sub_wire2(6, 75)    <= sub_wire11(75);
	sub_wire2(6, 76)    <= sub_wire11(76);
	sub_wire2(6, 77)    <= sub_wire11(77);
	sub_wire2(6, 78)    <= sub_wire11(78);
	sub_wire2(6, 79)    <= sub_wire11(79);
	sub_wire2(6, 80)    <= sub_wire11(80);
	sub_wire2(6, 81)    <= sub_wire11(81);
	sub_wire2(6, 82)    <= sub_wire11(82);
	sub_wire2(6, 83)    <= sub_wire11(83);
	sub_wire2(6, 84)    <= sub_wire11(84);
	sub_wire2(6, 85)    <= sub_wire11(85);
	sub_wire2(6, 86)    <= sub_wire11(86);
	sub_wire2(6, 87)    <= sub_wire11(87);
	sub_wire2(6, 88)    <= sub_wire11(88);
	sub_wire2(6, 89)    <= sub_wire11(89);
	sub_wire2(6, 90)    <= sub_wire11(90);
	sub_wire2(6, 91)    <= sub_wire11(91);
	sub_wire2(6, 92)    <= sub_wire11(92);
	sub_wire2(6, 93)    <= sub_wire11(93);
	sub_wire2(6, 94)    <= sub_wire11(94);
	sub_wire2(6, 95)    <= sub_wire11(95);
	sub_wire2(6, 96)    <= sub_wire11(96);
	sub_wire2(6, 97)    <= sub_wire11(97);
	sub_wire2(6, 98)    <= sub_wire11(98);
	sub_wire2(6, 99)    <= sub_wire11(99);
	sub_wire2(6, 100)    <= sub_wire11(100);
	sub_wire2(6, 101)    <= sub_wire11(101);
	sub_wire2(6, 102)    <= sub_wire11(102);
	sub_wire2(6, 103)    <= sub_wire11(103);
	sub_wire2(6, 104)    <= sub_wire11(104);
	sub_wire2(6, 105)    <= sub_wire11(105);
	sub_wire2(6, 106)    <= sub_wire11(106);
	sub_wire2(6, 107)    <= sub_wire11(107);
	sub_wire2(6, 108)    <= sub_wire11(108);
	sub_wire2(6, 109)    <= sub_wire11(109);
	sub_wire2(6, 110)    <= sub_wire11(110);
	sub_wire2(6, 111)    <= sub_wire11(111);
	sub_wire2(6, 112)    <= sub_wire11(112);
	sub_wire2(6, 113)    <= sub_wire11(113);
	sub_wire2(6, 114)    <= sub_wire11(114);
	sub_wire2(6, 115)    <= sub_wire11(115);
	sub_wire2(6, 116)    <= sub_wire11(116);
	sub_wire2(6, 117)    <= sub_wire11(117);
	sub_wire2(6, 118)    <= sub_wire11(118);
	sub_wire2(6, 119)    <= sub_wire11(119);
	sub_wire2(6, 120)    <= sub_wire11(120);
	sub_wire2(6, 121)    <= sub_wire11(121);
	sub_wire2(6, 122)    <= sub_wire11(122);
	sub_wire2(6, 123)    <= sub_wire11(123);
	sub_wire2(6, 124)    <= sub_wire11(124);
	sub_wire2(6, 125)    <= sub_wire11(125);
	sub_wire2(6, 126)    <= sub_wire11(126);
	sub_wire2(6, 127)    <= sub_wire11(127);
	sub_wire2(5, 0)    <= sub_wire12(0);
	sub_wire2(5, 1)    <= sub_wire12(1);
	sub_wire2(5, 2)    <= sub_wire12(2);
	sub_wire2(5, 3)    <= sub_wire12(3);
	sub_wire2(5, 4)    <= sub_wire12(4);
	sub_wire2(5, 5)    <= sub_wire12(5);
	sub_wire2(5, 6)    <= sub_wire12(6);
	sub_wire2(5, 7)    <= sub_wire12(7);
	sub_wire2(5, 8)    <= sub_wire12(8);
	sub_wire2(5, 9)    <= sub_wire12(9);
	sub_wire2(5, 10)    <= sub_wire12(10);
	sub_wire2(5, 11)    <= sub_wire12(11);
	sub_wire2(5, 12)    <= sub_wire12(12);
	sub_wire2(5, 13)    <= sub_wire12(13);
	sub_wire2(5, 14)    <= sub_wire12(14);
	sub_wire2(5, 15)    <= sub_wire12(15);
	sub_wire2(5, 16)    <= sub_wire12(16);
	sub_wire2(5, 17)    <= sub_wire12(17);
	sub_wire2(5, 18)    <= sub_wire12(18);
	sub_wire2(5, 19)    <= sub_wire12(19);
	sub_wire2(5, 20)    <= sub_wire12(20);
	sub_wire2(5, 21)    <= sub_wire12(21);
	sub_wire2(5, 22)    <= sub_wire12(22);
	sub_wire2(5, 23)    <= sub_wire12(23);
	sub_wire2(5, 24)    <= sub_wire12(24);
	sub_wire2(5, 25)    <= sub_wire12(25);
	sub_wire2(5, 26)    <= sub_wire12(26);
	sub_wire2(5, 27)    <= sub_wire12(27);
	sub_wire2(5, 28)    <= sub_wire12(28);
	sub_wire2(5, 29)    <= sub_wire12(29);
	sub_wire2(5, 30)    <= sub_wire12(30);
	sub_wire2(5, 31)    <= sub_wire12(31);
	sub_wire2(5, 32)    <= sub_wire12(32);
	sub_wire2(5, 33)    <= sub_wire12(33);
	sub_wire2(5, 34)    <= sub_wire12(34);
	sub_wire2(5, 35)    <= sub_wire12(35);
	sub_wire2(5, 36)    <= sub_wire12(36);
	sub_wire2(5, 37)    <= sub_wire12(37);
	sub_wire2(5, 38)    <= sub_wire12(38);
	sub_wire2(5, 39)    <= sub_wire12(39);
	sub_wire2(5, 40)    <= sub_wire12(40);
	sub_wire2(5, 41)    <= sub_wire12(41);
	sub_wire2(5, 42)    <= sub_wire12(42);
	sub_wire2(5, 43)    <= sub_wire12(43);
	sub_wire2(5, 44)    <= sub_wire12(44);
	sub_wire2(5, 45)    <= sub_wire12(45);
	sub_wire2(5, 46)    <= sub_wire12(46);
	sub_wire2(5, 47)    <= sub_wire12(47);
	sub_wire2(5, 48)    <= sub_wire12(48);
	sub_wire2(5, 49)    <= sub_wire12(49);
	sub_wire2(5, 50)    <= sub_wire12(50);
	sub_wire2(5, 51)    <= sub_wire12(51);
	sub_wire2(5, 52)    <= sub_wire12(52);
	sub_wire2(5, 53)    <= sub_wire12(53);
	sub_wire2(5, 54)    <= sub_wire12(54);
	sub_wire2(5, 55)    <= sub_wire12(55);
	sub_wire2(5, 56)    <= sub_wire12(56);
	sub_wire2(5, 57)    <= sub_wire12(57);
	sub_wire2(5, 58)    <= sub_wire12(58);
	sub_wire2(5, 59)    <= sub_wire12(59);
	sub_wire2(5, 60)    <= sub_wire12(60);
	sub_wire2(5, 61)    <= sub_wire12(61);
	sub_wire2(5, 62)    <= sub_wire12(62);
	sub_wire2(5, 63)    <= sub_wire12(63);
	sub_wire2(5, 64)    <= sub_wire12(64);
	sub_wire2(5, 65)    <= sub_wire12(65);
	sub_wire2(5, 66)    <= sub_wire12(66);
	sub_wire2(5, 67)    <= sub_wire12(67);
	sub_wire2(5, 68)    <= sub_wire12(68);
	sub_wire2(5, 69)    <= sub_wire12(69);
	sub_wire2(5, 70)    <= sub_wire12(70);
	sub_wire2(5, 71)    <= sub_wire12(71);
	sub_wire2(5, 72)    <= sub_wire12(72);
	sub_wire2(5, 73)    <= sub_wire12(73);
	sub_wire2(5, 74)    <= sub_wire12(74);
	sub_wire2(5, 75)    <= sub_wire12(75);
	sub_wire2(5, 76)    <= sub_wire12(76);
	sub_wire2(5, 77)    <= sub_wire12(77);
	sub_wire2(5, 78)    <= sub_wire12(78);
	sub_wire2(5, 79)    <= sub_wire12(79);
	sub_wire2(5, 80)    <= sub_wire12(80);
	sub_wire2(5, 81)    <= sub_wire12(81);
	sub_wire2(5, 82)    <= sub_wire12(82);
	sub_wire2(5, 83)    <= sub_wire12(83);
	sub_wire2(5, 84)    <= sub_wire12(84);
	sub_wire2(5, 85)    <= sub_wire12(85);
	sub_wire2(5, 86)    <= sub_wire12(86);
	sub_wire2(5, 87)    <= sub_wire12(87);
	sub_wire2(5, 88)    <= sub_wire12(88);
	sub_wire2(5, 89)    <= sub_wire12(89);
	sub_wire2(5, 90)    <= sub_wire12(90);
	sub_wire2(5, 91)    <= sub_wire12(91);
	sub_wire2(5, 92)    <= sub_wire12(92);
	sub_wire2(5, 93)    <= sub_wire12(93);
	sub_wire2(5, 94)    <= sub_wire12(94);
	sub_wire2(5, 95)    <= sub_wire12(95);
	sub_wire2(5, 96)    <= sub_wire12(96);
	sub_wire2(5, 97)    <= sub_wire12(97);
	sub_wire2(5, 98)    <= sub_wire12(98);
	sub_wire2(5, 99)    <= sub_wire12(99);
	sub_wire2(5, 100)    <= sub_wire12(100);
	sub_wire2(5, 101)    <= sub_wire12(101);
	sub_wire2(5, 102)    <= sub_wire12(102);
	sub_wire2(5, 103)    <= sub_wire12(103);
	sub_wire2(5, 104)    <= sub_wire12(104);
	sub_wire2(5, 105)    <= sub_wire12(105);
	sub_wire2(5, 106)    <= sub_wire12(106);
	sub_wire2(5, 107)    <= sub_wire12(107);
	sub_wire2(5, 108)    <= sub_wire12(108);
	sub_wire2(5, 109)    <= sub_wire12(109);
	sub_wire2(5, 110)    <= sub_wire12(110);
	sub_wire2(5, 111)    <= sub_wire12(111);
	sub_wire2(5, 112)    <= sub_wire12(112);
	sub_wire2(5, 113)    <= sub_wire12(113);
	sub_wire2(5, 114)    <= sub_wire12(114);
	sub_wire2(5, 115)    <= sub_wire12(115);
	sub_wire2(5, 116)    <= sub_wire12(116);
	sub_wire2(5, 117)    <= sub_wire12(117);
	sub_wire2(5, 118)    <= sub_wire12(118);
	sub_wire2(5, 119)    <= sub_wire12(119);
	sub_wire2(5, 120)    <= sub_wire12(120);
	sub_wire2(5, 121)    <= sub_wire12(121);
	sub_wire2(5, 122)    <= sub_wire12(122);
	sub_wire2(5, 123)    <= sub_wire12(123);
	sub_wire2(5, 124)    <= sub_wire12(124);
	sub_wire2(5, 125)    <= sub_wire12(125);
	sub_wire2(5, 126)    <= sub_wire12(126);
	sub_wire2(5, 127)    <= sub_wire12(127);
	sub_wire2(4, 0)    <= sub_wire13(0);
	sub_wire2(4, 1)    <= sub_wire13(1);
	sub_wire2(4, 2)    <= sub_wire13(2);
	sub_wire2(4, 3)    <= sub_wire13(3);
	sub_wire2(4, 4)    <= sub_wire13(4);
	sub_wire2(4, 5)    <= sub_wire13(5);
	sub_wire2(4, 6)    <= sub_wire13(6);
	sub_wire2(4, 7)    <= sub_wire13(7);
	sub_wire2(4, 8)    <= sub_wire13(8);
	sub_wire2(4, 9)    <= sub_wire13(9);
	sub_wire2(4, 10)    <= sub_wire13(10);
	sub_wire2(4, 11)    <= sub_wire13(11);
	sub_wire2(4, 12)    <= sub_wire13(12);
	sub_wire2(4, 13)    <= sub_wire13(13);
	sub_wire2(4, 14)    <= sub_wire13(14);
	sub_wire2(4, 15)    <= sub_wire13(15);
	sub_wire2(4, 16)    <= sub_wire13(16);
	sub_wire2(4, 17)    <= sub_wire13(17);
	sub_wire2(4, 18)    <= sub_wire13(18);
	sub_wire2(4, 19)    <= sub_wire13(19);
	sub_wire2(4, 20)    <= sub_wire13(20);
	sub_wire2(4, 21)    <= sub_wire13(21);
	sub_wire2(4, 22)    <= sub_wire13(22);
	sub_wire2(4, 23)    <= sub_wire13(23);
	sub_wire2(4, 24)    <= sub_wire13(24);
	sub_wire2(4, 25)    <= sub_wire13(25);
	sub_wire2(4, 26)    <= sub_wire13(26);
	sub_wire2(4, 27)    <= sub_wire13(27);
	sub_wire2(4, 28)    <= sub_wire13(28);
	sub_wire2(4, 29)    <= sub_wire13(29);
	sub_wire2(4, 30)    <= sub_wire13(30);
	sub_wire2(4, 31)    <= sub_wire13(31);
	sub_wire2(4, 32)    <= sub_wire13(32);
	sub_wire2(4, 33)    <= sub_wire13(33);
	sub_wire2(4, 34)    <= sub_wire13(34);
	sub_wire2(4, 35)    <= sub_wire13(35);
	sub_wire2(4, 36)    <= sub_wire13(36);
	sub_wire2(4, 37)    <= sub_wire13(37);
	sub_wire2(4, 38)    <= sub_wire13(38);
	sub_wire2(4, 39)    <= sub_wire13(39);
	sub_wire2(4, 40)    <= sub_wire13(40);
	sub_wire2(4, 41)    <= sub_wire13(41);
	sub_wire2(4, 42)    <= sub_wire13(42);
	sub_wire2(4, 43)    <= sub_wire13(43);
	sub_wire2(4, 44)    <= sub_wire13(44);
	sub_wire2(4, 45)    <= sub_wire13(45);
	sub_wire2(4, 46)    <= sub_wire13(46);
	sub_wire2(4, 47)    <= sub_wire13(47);
	sub_wire2(4, 48)    <= sub_wire13(48);
	sub_wire2(4, 49)    <= sub_wire13(49);
	sub_wire2(4, 50)    <= sub_wire13(50);
	sub_wire2(4, 51)    <= sub_wire13(51);
	sub_wire2(4, 52)    <= sub_wire13(52);
	sub_wire2(4, 53)    <= sub_wire13(53);
	sub_wire2(4, 54)    <= sub_wire13(54);
	sub_wire2(4, 55)    <= sub_wire13(55);
	sub_wire2(4, 56)    <= sub_wire13(56);
	sub_wire2(4, 57)    <= sub_wire13(57);
	sub_wire2(4, 58)    <= sub_wire13(58);
	sub_wire2(4, 59)    <= sub_wire13(59);
	sub_wire2(4, 60)    <= sub_wire13(60);
	sub_wire2(4, 61)    <= sub_wire13(61);
	sub_wire2(4, 62)    <= sub_wire13(62);
	sub_wire2(4, 63)    <= sub_wire13(63);
	sub_wire2(4, 64)    <= sub_wire13(64);
	sub_wire2(4, 65)    <= sub_wire13(65);
	sub_wire2(4, 66)    <= sub_wire13(66);
	sub_wire2(4, 67)    <= sub_wire13(67);
	sub_wire2(4, 68)    <= sub_wire13(68);
	sub_wire2(4, 69)    <= sub_wire13(69);
	sub_wire2(4, 70)    <= sub_wire13(70);
	sub_wire2(4, 71)    <= sub_wire13(71);
	sub_wire2(4, 72)    <= sub_wire13(72);
	sub_wire2(4, 73)    <= sub_wire13(73);
	sub_wire2(4, 74)    <= sub_wire13(74);
	sub_wire2(4, 75)    <= sub_wire13(75);
	sub_wire2(4, 76)    <= sub_wire13(76);
	sub_wire2(4, 77)    <= sub_wire13(77);
	sub_wire2(4, 78)    <= sub_wire13(78);
	sub_wire2(4, 79)    <= sub_wire13(79);
	sub_wire2(4, 80)    <= sub_wire13(80);
	sub_wire2(4, 81)    <= sub_wire13(81);
	sub_wire2(4, 82)    <= sub_wire13(82);
	sub_wire2(4, 83)    <= sub_wire13(83);
	sub_wire2(4, 84)    <= sub_wire13(84);
	sub_wire2(4, 85)    <= sub_wire13(85);
	sub_wire2(4, 86)    <= sub_wire13(86);
	sub_wire2(4, 87)    <= sub_wire13(87);
	sub_wire2(4, 88)    <= sub_wire13(88);
	sub_wire2(4, 89)    <= sub_wire13(89);
	sub_wire2(4, 90)    <= sub_wire13(90);
	sub_wire2(4, 91)    <= sub_wire13(91);
	sub_wire2(4, 92)    <= sub_wire13(92);
	sub_wire2(4, 93)    <= sub_wire13(93);
	sub_wire2(4, 94)    <= sub_wire13(94);
	sub_wire2(4, 95)    <= sub_wire13(95);
	sub_wire2(4, 96)    <= sub_wire13(96);
	sub_wire2(4, 97)    <= sub_wire13(97);
	sub_wire2(4, 98)    <= sub_wire13(98);
	sub_wire2(4, 99)    <= sub_wire13(99);
	sub_wire2(4, 100)    <= sub_wire13(100);
	sub_wire2(4, 101)    <= sub_wire13(101);
	sub_wire2(4, 102)    <= sub_wire13(102);
	sub_wire2(4, 103)    <= sub_wire13(103);
	sub_wire2(4, 104)    <= sub_wire13(104);
	sub_wire2(4, 105)    <= sub_wire13(105);
	sub_wire2(4, 106)    <= sub_wire13(106);
	sub_wire2(4, 107)    <= sub_wire13(107);
	sub_wire2(4, 108)    <= sub_wire13(108);
	sub_wire2(4, 109)    <= sub_wire13(109);
	sub_wire2(4, 110)    <= sub_wire13(110);
	sub_wire2(4, 111)    <= sub_wire13(111);
	sub_wire2(4, 112)    <= sub_wire13(112);
	sub_wire2(4, 113)    <= sub_wire13(113);
	sub_wire2(4, 114)    <= sub_wire13(114);
	sub_wire2(4, 115)    <= sub_wire13(115);
	sub_wire2(4, 116)    <= sub_wire13(116);
	sub_wire2(4, 117)    <= sub_wire13(117);
	sub_wire2(4, 118)    <= sub_wire13(118);
	sub_wire2(4, 119)    <= sub_wire13(119);
	sub_wire2(4, 120)    <= sub_wire13(120);
	sub_wire2(4, 121)    <= sub_wire13(121);
	sub_wire2(4, 122)    <= sub_wire13(122);
	sub_wire2(4, 123)    <= sub_wire13(123);
	sub_wire2(4, 124)    <= sub_wire13(124);
	sub_wire2(4, 125)    <= sub_wire13(125);
	sub_wire2(4, 126)    <= sub_wire13(126);
	sub_wire2(4, 127)    <= sub_wire13(127);
	sub_wire2(3, 0)    <= sub_wire14(0);
	sub_wire2(3, 1)    <= sub_wire14(1);
	sub_wire2(3, 2)    <= sub_wire14(2);
	sub_wire2(3, 3)    <= sub_wire14(3);
	sub_wire2(3, 4)    <= sub_wire14(4);
	sub_wire2(3, 5)    <= sub_wire14(5);
	sub_wire2(3, 6)    <= sub_wire14(6);
	sub_wire2(3, 7)    <= sub_wire14(7);
	sub_wire2(3, 8)    <= sub_wire14(8);
	sub_wire2(3, 9)    <= sub_wire14(9);
	sub_wire2(3, 10)    <= sub_wire14(10);
	sub_wire2(3, 11)    <= sub_wire14(11);
	sub_wire2(3, 12)    <= sub_wire14(12);
	sub_wire2(3, 13)    <= sub_wire14(13);
	sub_wire2(3, 14)    <= sub_wire14(14);
	sub_wire2(3, 15)    <= sub_wire14(15);
	sub_wire2(3, 16)    <= sub_wire14(16);
	sub_wire2(3, 17)    <= sub_wire14(17);
	sub_wire2(3, 18)    <= sub_wire14(18);
	sub_wire2(3, 19)    <= sub_wire14(19);
	sub_wire2(3, 20)    <= sub_wire14(20);
	sub_wire2(3, 21)    <= sub_wire14(21);
	sub_wire2(3, 22)    <= sub_wire14(22);
	sub_wire2(3, 23)    <= sub_wire14(23);
	sub_wire2(3, 24)    <= sub_wire14(24);
	sub_wire2(3, 25)    <= sub_wire14(25);
	sub_wire2(3, 26)    <= sub_wire14(26);
	sub_wire2(3, 27)    <= sub_wire14(27);
	sub_wire2(3, 28)    <= sub_wire14(28);
	sub_wire2(3, 29)    <= sub_wire14(29);
	sub_wire2(3, 30)    <= sub_wire14(30);
	sub_wire2(3, 31)    <= sub_wire14(31);
	sub_wire2(3, 32)    <= sub_wire14(32);
	sub_wire2(3, 33)    <= sub_wire14(33);
	sub_wire2(3, 34)    <= sub_wire14(34);
	sub_wire2(3, 35)    <= sub_wire14(35);
	sub_wire2(3, 36)    <= sub_wire14(36);
	sub_wire2(3, 37)    <= sub_wire14(37);
	sub_wire2(3, 38)    <= sub_wire14(38);
	sub_wire2(3, 39)    <= sub_wire14(39);
	sub_wire2(3, 40)    <= sub_wire14(40);
	sub_wire2(3, 41)    <= sub_wire14(41);
	sub_wire2(3, 42)    <= sub_wire14(42);
	sub_wire2(3, 43)    <= sub_wire14(43);
	sub_wire2(3, 44)    <= sub_wire14(44);
	sub_wire2(3, 45)    <= sub_wire14(45);
	sub_wire2(3, 46)    <= sub_wire14(46);
	sub_wire2(3, 47)    <= sub_wire14(47);
	sub_wire2(3, 48)    <= sub_wire14(48);
	sub_wire2(3, 49)    <= sub_wire14(49);
	sub_wire2(3, 50)    <= sub_wire14(50);
	sub_wire2(3, 51)    <= sub_wire14(51);
	sub_wire2(3, 52)    <= sub_wire14(52);
	sub_wire2(3, 53)    <= sub_wire14(53);
	sub_wire2(3, 54)    <= sub_wire14(54);
	sub_wire2(3, 55)    <= sub_wire14(55);
	sub_wire2(3, 56)    <= sub_wire14(56);
	sub_wire2(3, 57)    <= sub_wire14(57);
	sub_wire2(3, 58)    <= sub_wire14(58);
	sub_wire2(3, 59)    <= sub_wire14(59);
	sub_wire2(3, 60)    <= sub_wire14(60);
	sub_wire2(3, 61)    <= sub_wire14(61);
	sub_wire2(3, 62)    <= sub_wire14(62);
	sub_wire2(3, 63)    <= sub_wire14(63);
	sub_wire2(3, 64)    <= sub_wire14(64);
	sub_wire2(3, 65)    <= sub_wire14(65);
	sub_wire2(3, 66)    <= sub_wire14(66);
	sub_wire2(3, 67)    <= sub_wire14(67);
	sub_wire2(3, 68)    <= sub_wire14(68);
	sub_wire2(3, 69)    <= sub_wire14(69);
	sub_wire2(3, 70)    <= sub_wire14(70);
	sub_wire2(3, 71)    <= sub_wire14(71);
	sub_wire2(3, 72)    <= sub_wire14(72);
	sub_wire2(3, 73)    <= sub_wire14(73);
	sub_wire2(3, 74)    <= sub_wire14(74);
	sub_wire2(3, 75)    <= sub_wire14(75);
	sub_wire2(3, 76)    <= sub_wire14(76);
	sub_wire2(3, 77)    <= sub_wire14(77);
	sub_wire2(3, 78)    <= sub_wire14(78);
	sub_wire2(3, 79)    <= sub_wire14(79);
	sub_wire2(3, 80)    <= sub_wire14(80);
	sub_wire2(3, 81)    <= sub_wire14(81);
	sub_wire2(3, 82)    <= sub_wire14(82);
	sub_wire2(3, 83)    <= sub_wire14(83);
	sub_wire2(3, 84)    <= sub_wire14(84);
	sub_wire2(3, 85)    <= sub_wire14(85);
	sub_wire2(3, 86)    <= sub_wire14(86);
	sub_wire2(3, 87)    <= sub_wire14(87);
	sub_wire2(3, 88)    <= sub_wire14(88);
	sub_wire2(3, 89)    <= sub_wire14(89);
	sub_wire2(3, 90)    <= sub_wire14(90);
	sub_wire2(3, 91)    <= sub_wire14(91);
	sub_wire2(3, 92)    <= sub_wire14(92);
	sub_wire2(3, 93)    <= sub_wire14(93);
	sub_wire2(3, 94)    <= sub_wire14(94);
	sub_wire2(3, 95)    <= sub_wire14(95);
	sub_wire2(3, 96)    <= sub_wire14(96);
	sub_wire2(3, 97)    <= sub_wire14(97);
	sub_wire2(3, 98)    <= sub_wire14(98);
	sub_wire2(3, 99)    <= sub_wire14(99);
	sub_wire2(3, 100)    <= sub_wire14(100);
	sub_wire2(3, 101)    <= sub_wire14(101);
	sub_wire2(3, 102)    <= sub_wire14(102);
	sub_wire2(3, 103)    <= sub_wire14(103);
	sub_wire2(3, 104)    <= sub_wire14(104);
	sub_wire2(3, 105)    <= sub_wire14(105);
	sub_wire2(3, 106)    <= sub_wire14(106);
	sub_wire2(3, 107)    <= sub_wire14(107);
	sub_wire2(3, 108)    <= sub_wire14(108);
	sub_wire2(3, 109)    <= sub_wire14(109);
	sub_wire2(3, 110)    <= sub_wire14(110);
	sub_wire2(3, 111)    <= sub_wire14(111);
	sub_wire2(3, 112)    <= sub_wire14(112);
	sub_wire2(3, 113)    <= sub_wire14(113);
	sub_wire2(3, 114)    <= sub_wire14(114);
	sub_wire2(3, 115)    <= sub_wire14(115);
	sub_wire2(3, 116)    <= sub_wire14(116);
	sub_wire2(3, 117)    <= sub_wire14(117);
	sub_wire2(3, 118)    <= sub_wire14(118);
	sub_wire2(3, 119)    <= sub_wire14(119);
	sub_wire2(3, 120)    <= sub_wire14(120);
	sub_wire2(3, 121)    <= sub_wire14(121);
	sub_wire2(3, 122)    <= sub_wire14(122);
	sub_wire2(3, 123)    <= sub_wire14(123);
	sub_wire2(3, 124)    <= sub_wire14(124);
	sub_wire2(3, 125)    <= sub_wire14(125);
	sub_wire2(3, 126)    <= sub_wire14(126);
	sub_wire2(3, 127)    <= sub_wire14(127);
	sub_wire2(2, 0)    <= sub_wire15(0);
	sub_wire2(2, 1)    <= sub_wire15(1);
	sub_wire2(2, 2)    <= sub_wire15(2);
	sub_wire2(2, 3)    <= sub_wire15(3);
	sub_wire2(2, 4)    <= sub_wire15(4);
	sub_wire2(2, 5)    <= sub_wire15(5);
	sub_wire2(2, 6)    <= sub_wire15(6);
	sub_wire2(2, 7)    <= sub_wire15(7);
	sub_wire2(2, 8)    <= sub_wire15(8);
	sub_wire2(2, 9)    <= sub_wire15(9);
	sub_wire2(2, 10)    <= sub_wire15(10);
	sub_wire2(2, 11)    <= sub_wire15(11);
	sub_wire2(2, 12)    <= sub_wire15(12);
	sub_wire2(2, 13)    <= sub_wire15(13);
	sub_wire2(2, 14)    <= sub_wire15(14);
	sub_wire2(2, 15)    <= sub_wire15(15);
	sub_wire2(2, 16)    <= sub_wire15(16);
	sub_wire2(2, 17)    <= sub_wire15(17);
	sub_wire2(2, 18)    <= sub_wire15(18);
	sub_wire2(2, 19)    <= sub_wire15(19);
	sub_wire2(2, 20)    <= sub_wire15(20);
	sub_wire2(2, 21)    <= sub_wire15(21);
	sub_wire2(2, 22)    <= sub_wire15(22);
	sub_wire2(2, 23)    <= sub_wire15(23);
	sub_wire2(2, 24)    <= sub_wire15(24);
	sub_wire2(2, 25)    <= sub_wire15(25);
	sub_wire2(2, 26)    <= sub_wire15(26);
	sub_wire2(2, 27)    <= sub_wire15(27);
	sub_wire2(2, 28)    <= sub_wire15(28);
	sub_wire2(2, 29)    <= sub_wire15(29);
	sub_wire2(2, 30)    <= sub_wire15(30);
	sub_wire2(2, 31)    <= sub_wire15(31);
	sub_wire2(2, 32)    <= sub_wire15(32);
	sub_wire2(2, 33)    <= sub_wire15(33);
	sub_wire2(2, 34)    <= sub_wire15(34);
	sub_wire2(2, 35)    <= sub_wire15(35);
	sub_wire2(2, 36)    <= sub_wire15(36);
	sub_wire2(2, 37)    <= sub_wire15(37);
	sub_wire2(2, 38)    <= sub_wire15(38);
	sub_wire2(2, 39)    <= sub_wire15(39);
	sub_wire2(2, 40)    <= sub_wire15(40);
	sub_wire2(2, 41)    <= sub_wire15(41);
	sub_wire2(2, 42)    <= sub_wire15(42);
	sub_wire2(2, 43)    <= sub_wire15(43);
	sub_wire2(2, 44)    <= sub_wire15(44);
	sub_wire2(2, 45)    <= sub_wire15(45);
	sub_wire2(2, 46)    <= sub_wire15(46);
	sub_wire2(2, 47)    <= sub_wire15(47);
	sub_wire2(2, 48)    <= sub_wire15(48);
	sub_wire2(2, 49)    <= sub_wire15(49);
	sub_wire2(2, 50)    <= sub_wire15(50);
	sub_wire2(2, 51)    <= sub_wire15(51);
	sub_wire2(2, 52)    <= sub_wire15(52);
	sub_wire2(2, 53)    <= sub_wire15(53);
	sub_wire2(2, 54)    <= sub_wire15(54);
	sub_wire2(2, 55)    <= sub_wire15(55);
	sub_wire2(2, 56)    <= sub_wire15(56);
	sub_wire2(2, 57)    <= sub_wire15(57);
	sub_wire2(2, 58)    <= sub_wire15(58);
	sub_wire2(2, 59)    <= sub_wire15(59);
	sub_wire2(2, 60)    <= sub_wire15(60);
	sub_wire2(2, 61)    <= sub_wire15(61);
	sub_wire2(2, 62)    <= sub_wire15(62);
	sub_wire2(2, 63)    <= sub_wire15(63);
	sub_wire2(2, 64)    <= sub_wire15(64);
	sub_wire2(2, 65)    <= sub_wire15(65);
	sub_wire2(2, 66)    <= sub_wire15(66);
	sub_wire2(2, 67)    <= sub_wire15(67);
	sub_wire2(2, 68)    <= sub_wire15(68);
	sub_wire2(2, 69)    <= sub_wire15(69);
	sub_wire2(2, 70)    <= sub_wire15(70);
	sub_wire2(2, 71)    <= sub_wire15(71);
	sub_wire2(2, 72)    <= sub_wire15(72);
	sub_wire2(2, 73)    <= sub_wire15(73);
	sub_wire2(2, 74)    <= sub_wire15(74);
	sub_wire2(2, 75)    <= sub_wire15(75);
	sub_wire2(2, 76)    <= sub_wire15(76);
	sub_wire2(2, 77)    <= sub_wire15(77);
	sub_wire2(2, 78)    <= sub_wire15(78);
	sub_wire2(2, 79)    <= sub_wire15(79);
	sub_wire2(2, 80)    <= sub_wire15(80);
	sub_wire2(2, 81)    <= sub_wire15(81);
	sub_wire2(2, 82)    <= sub_wire15(82);
	sub_wire2(2, 83)    <= sub_wire15(83);
	sub_wire2(2, 84)    <= sub_wire15(84);
	sub_wire2(2, 85)    <= sub_wire15(85);
	sub_wire2(2, 86)    <= sub_wire15(86);
	sub_wire2(2, 87)    <= sub_wire15(87);
	sub_wire2(2, 88)    <= sub_wire15(88);
	sub_wire2(2, 89)    <= sub_wire15(89);
	sub_wire2(2, 90)    <= sub_wire15(90);
	sub_wire2(2, 91)    <= sub_wire15(91);
	sub_wire2(2, 92)    <= sub_wire15(92);
	sub_wire2(2, 93)    <= sub_wire15(93);
	sub_wire2(2, 94)    <= sub_wire15(94);
	sub_wire2(2, 95)    <= sub_wire15(95);
	sub_wire2(2, 96)    <= sub_wire15(96);
	sub_wire2(2, 97)    <= sub_wire15(97);
	sub_wire2(2, 98)    <= sub_wire15(98);
	sub_wire2(2, 99)    <= sub_wire15(99);
	sub_wire2(2, 100)    <= sub_wire15(100);
	sub_wire2(2, 101)    <= sub_wire15(101);
	sub_wire2(2, 102)    <= sub_wire15(102);
	sub_wire2(2, 103)    <= sub_wire15(103);
	sub_wire2(2, 104)    <= sub_wire15(104);
	sub_wire2(2, 105)    <= sub_wire15(105);
	sub_wire2(2, 106)    <= sub_wire15(106);
	sub_wire2(2, 107)    <= sub_wire15(107);
	sub_wire2(2, 108)    <= sub_wire15(108);
	sub_wire2(2, 109)    <= sub_wire15(109);
	sub_wire2(2, 110)    <= sub_wire15(110);
	sub_wire2(2, 111)    <= sub_wire15(111);
	sub_wire2(2, 112)    <= sub_wire15(112);
	sub_wire2(2, 113)    <= sub_wire15(113);
	sub_wire2(2, 114)    <= sub_wire15(114);
	sub_wire2(2, 115)    <= sub_wire15(115);
	sub_wire2(2, 116)    <= sub_wire15(116);
	sub_wire2(2, 117)    <= sub_wire15(117);
	sub_wire2(2, 118)    <= sub_wire15(118);
	sub_wire2(2, 119)    <= sub_wire15(119);
	sub_wire2(2, 120)    <= sub_wire15(120);
	sub_wire2(2, 121)    <= sub_wire15(121);
	sub_wire2(2, 122)    <= sub_wire15(122);
	sub_wire2(2, 123)    <= sub_wire15(123);
	sub_wire2(2, 124)    <= sub_wire15(124);
	sub_wire2(2, 125)    <= sub_wire15(125);
	sub_wire2(2, 126)    <= sub_wire15(126);
	sub_wire2(2, 127)    <= sub_wire15(127);
	sub_wire2(1, 0)    <= sub_wire16(0);
	sub_wire2(1, 1)    <= sub_wire16(1);
	sub_wire2(1, 2)    <= sub_wire16(2);
	sub_wire2(1, 3)    <= sub_wire16(3);
	sub_wire2(1, 4)    <= sub_wire16(4);
	sub_wire2(1, 5)    <= sub_wire16(5);
	sub_wire2(1, 6)    <= sub_wire16(6);
	sub_wire2(1, 7)    <= sub_wire16(7);
	sub_wire2(1, 8)    <= sub_wire16(8);
	sub_wire2(1, 9)    <= sub_wire16(9);
	sub_wire2(1, 10)    <= sub_wire16(10);
	sub_wire2(1, 11)    <= sub_wire16(11);
	sub_wire2(1, 12)    <= sub_wire16(12);
	sub_wire2(1, 13)    <= sub_wire16(13);
	sub_wire2(1, 14)    <= sub_wire16(14);
	sub_wire2(1, 15)    <= sub_wire16(15);
	sub_wire2(1, 16)    <= sub_wire16(16);
	sub_wire2(1, 17)    <= sub_wire16(17);
	sub_wire2(1, 18)    <= sub_wire16(18);
	sub_wire2(1, 19)    <= sub_wire16(19);
	sub_wire2(1, 20)    <= sub_wire16(20);
	sub_wire2(1, 21)    <= sub_wire16(21);
	sub_wire2(1, 22)    <= sub_wire16(22);
	sub_wire2(1, 23)    <= sub_wire16(23);
	sub_wire2(1, 24)    <= sub_wire16(24);
	sub_wire2(1, 25)    <= sub_wire16(25);
	sub_wire2(1, 26)    <= sub_wire16(26);
	sub_wire2(1, 27)    <= sub_wire16(27);
	sub_wire2(1, 28)    <= sub_wire16(28);
	sub_wire2(1, 29)    <= sub_wire16(29);
	sub_wire2(1, 30)    <= sub_wire16(30);
	sub_wire2(1, 31)    <= sub_wire16(31);
	sub_wire2(1, 32)    <= sub_wire16(32);
	sub_wire2(1, 33)    <= sub_wire16(33);
	sub_wire2(1, 34)    <= sub_wire16(34);
	sub_wire2(1, 35)    <= sub_wire16(35);
	sub_wire2(1, 36)    <= sub_wire16(36);
	sub_wire2(1, 37)    <= sub_wire16(37);
	sub_wire2(1, 38)    <= sub_wire16(38);
	sub_wire2(1, 39)    <= sub_wire16(39);
	sub_wire2(1, 40)    <= sub_wire16(40);
	sub_wire2(1, 41)    <= sub_wire16(41);
	sub_wire2(1, 42)    <= sub_wire16(42);
	sub_wire2(1, 43)    <= sub_wire16(43);
	sub_wire2(1, 44)    <= sub_wire16(44);
	sub_wire2(1, 45)    <= sub_wire16(45);
	sub_wire2(1, 46)    <= sub_wire16(46);
	sub_wire2(1, 47)    <= sub_wire16(47);
	sub_wire2(1, 48)    <= sub_wire16(48);
	sub_wire2(1, 49)    <= sub_wire16(49);
	sub_wire2(1, 50)    <= sub_wire16(50);
	sub_wire2(1, 51)    <= sub_wire16(51);
	sub_wire2(1, 52)    <= sub_wire16(52);
	sub_wire2(1, 53)    <= sub_wire16(53);
	sub_wire2(1, 54)    <= sub_wire16(54);
	sub_wire2(1, 55)    <= sub_wire16(55);
	sub_wire2(1, 56)    <= sub_wire16(56);
	sub_wire2(1, 57)    <= sub_wire16(57);
	sub_wire2(1, 58)    <= sub_wire16(58);
	sub_wire2(1, 59)    <= sub_wire16(59);
	sub_wire2(1, 60)    <= sub_wire16(60);
	sub_wire2(1, 61)    <= sub_wire16(61);
	sub_wire2(1, 62)    <= sub_wire16(62);
	sub_wire2(1, 63)    <= sub_wire16(63);
	sub_wire2(1, 64)    <= sub_wire16(64);
	sub_wire2(1, 65)    <= sub_wire16(65);
	sub_wire2(1, 66)    <= sub_wire16(66);
	sub_wire2(1, 67)    <= sub_wire16(67);
	sub_wire2(1, 68)    <= sub_wire16(68);
	sub_wire2(1, 69)    <= sub_wire16(69);
	sub_wire2(1, 70)    <= sub_wire16(70);
	sub_wire2(1, 71)    <= sub_wire16(71);
	sub_wire2(1, 72)    <= sub_wire16(72);
	sub_wire2(1, 73)    <= sub_wire16(73);
	sub_wire2(1, 74)    <= sub_wire16(74);
	sub_wire2(1, 75)    <= sub_wire16(75);
	sub_wire2(1, 76)    <= sub_wire16(76);
	sub_wire2(1, 77)    <= sub_wire16(77);
	sub_wire2(1, 78)    <= sub_wire16(78);
	sub_wire2(1, 79)    <= sub_wire16(79);
	sub_wire2(1, 80)    <= sub_wire16(80);
	sub_wire2(1, 81)    <= sub_wire16(81);
	sub_wire2(1, 82)    <= sub_wire16(82);
	sub_wire2(1, 83)    <= sub_wire16(83);
	sub_wire2(1, 84)    <= sub_wire16(84);
	sub_wire2(1, 85)    <= sub_wire16(85);
	sub_wire2(1, 86)    <= sub_wire16(86);
	sub_wire2(1, 87)    <= sub_wire16(87);
	sub_wire2(1, 88)    <= sub_wire16(88);
	sub_wire2(1, 89)    <= sub_wire16(89);
	sub_wire2(1, 90)    <= sub_wire16(90);
	sub_wire2(1, 91)    <= sub_wire16(91);
	sub_wire2(1, 92)    <= sub_wire16(92);
	sub_wire2(1, 93)    <= sub_wire16(93);
	sub_wire2(1, 94)    <= sub_wire16(94);
	sub_wire2(1, 95)    <= sub_wire16(95);
	sub_wire2(1, 96)    <= sub_wire16(96);
	sub_wire2(1, 97)    <= sub_wire16(97);
	sub_wire2(1, 98)    <= sub_wire16(98);
	sub_wire2(1, 99)    <= sub_wire16(99);
	sub_wire2(1, 100)    <= sub_wire16(100);
	sub_wire2(1, 101)    <= sub_wire16(101);
	sub_wire2(1, 102)    <= sub_wire16(102);
	sub_wire2(1, 103)    <= sub_wire16(103);
	sub_wire2(1, 104)    <= sub_wire16(104);
	sub_wire2(1, 105)    <= sub_wire16(105);
	sub_wire2(1, 106)    <= sub_wire16(106);
	sub_wire2(1, 107)    <= sub_wire16(107);
	sub_wire2(1, 108)    <= sub_wire16(108);
	sub_wire2(1, 109)    <= sub_wire16(109);
	sub_wire2(1, 110)    <= sub_wire16(110);
	sub_wire2(1, 111)    <= sub_wire16(111);
	sub_wire2(1, 112)    <= sub_wire16(112);
	sub_wire2(1, 113)    <= sub_wire16(113);
	sub_wire2(1, 114)    <= sub_wire16(114);
	sub_wire2(1, 115)    <= sub_wire16(115);
	sub_wire2(1, 116)    <= sub_wire16(116);
	sub_wire2(1, 117)    <= sub_wire16(117);
	sub_wire2(1, 118)    <= sub_wire16(118);
	sub_wire2(1, 119)    <= sub_wire16(119);
	sub_wire2(1, 120)    <= sub_wire16(120);
	sub_wire2(1, 121)    <= sub_wire16(121);
	sub_wire2(1, 122)    <= sub_wire16(122);
	sub_wire2(1, 123)    <= sub_wire16(123);
	sub_wire2(1, 124)    <= sub_wire16(124);
	sub_wire2(1, 125)    <= sub_wire16(125);
	sub_wire2(1, 126)    <= sub_wire16(126);
	sub_wire2(1, 127)    <= sub_wire16(127);
	sub_wire2(0, 0)    <= sub_wire17(0);
	sub_wire2(0, 1)    <= sub_wire17(1);
	sub_wire2(0, 2)    <= sub_wire17(2);
	sub_wire2(0, 3)    <= sub_wire17(3);
	sub_wire2(0, 4)    <= sub_wire17(4);
	sub_wire2(0, 5)    <= sub_wire17(5);
	sub_wire2(0, 6)    <= sub_wire17(6);
	sub_wire2(0, 7)    <= sub_wire17(7);
	sub_wire2(0, 8)    <= sub_wire17(8);
	sub_wire2(0, 9)    <= sub_wire17(9);
	sub_wire2(0, 10)    <= sub_wire17(10);
	sub_wire2(0, 11)    <= sub_wire17(11);
	sub_wire2(0, 12)    <= sub_wire17(12);
	sub_wire2(0, 13)    <= sub_wire17(13);
	sub_wire2(0, 14)    <= sub_wire17(14);
	sub_wire2(0, 15)    <= sub_wire17(15);
	sub_wire2(0, 16)    <= sub_wire17(16);
	sub_wire2(0, 17)    <= sub_wire17(17);
	sub_wire2(0, 18)    <= sub_wire17(18);
	sub_wire2(0, 19)    <= sub_wire17(19);
	sub_wire2(0, 20)    <= sub_wire17(20);
	sub_wire2(0, 21)    <= sub_wire17(21);
	sub_wire2(0, 22)    <= sub_wire17(22);
	sub_wire2(0, 23)    <= sub_wire17(23);
	sub_wire2(0, 24)    <= sub_wire17(24);
	sub_wire2(0, 25)    <= sub_wire17(25);
	sub_wire2(0, 26)    <= sub_wire17(26);
	sub_wire2(0, 27)    <= sub_wire17(27);
	sub_wire2(0, 28)    <= sub_wire17(28);
	sub_wire2(0, 29)    <= sub_wire17(29);
	sub_wire2(0, 30)    <= sub_wire17(30);
	sub_wire2(0, 31)    <= sub_wire17(31);
	sub_wire2(0, 32)    <= sub_wire17(32);
	sub_wire2(0, 33)    <= sub_wire17(33);
	sub_wire2(0, 34)    <= sub_wire17(34);
	sub_wire2(0, 35)    <= sub_wire17(35);
	sub_wire2(0, 36)    <= sub_wire17(36);
	sub_wire2(0, 37)    <= sub_wire17(37);
	sub_wire2(0, 38)    <= sub_wire17(38);
	sub_wire2(0, 39)    <= sub_wire17(39);
	sub_wire2(0, 40)    <= sub_wire17(40);
	sub_wire2(0, 41)    <= sub_wire17(41);
	sub_wire2(0, 42)    <= sub_wire17(42);
	sub_wire2(0, 43)    <= sub_wire17(43);
	sub_wire2(0, 44)    <= sub_wire17(44);
	sub_wire2(0, 45)    <= sub_wire17(45);
	sub_wire2(0, 46)    <= sub_wire17(46);
	sub_wire2(0, 47)    <= sub_wire17(47);
	sub_wire2(0, 48)    <= sub_wire17(48);
	sub_wire2(0, 49)    <= sub_wire17(49);
	sub_wire2(0, 50)    <= sub_wire17(50);
	sub_wire2(0, 51)    <= sub_wire17(51);
	sub_wire2(0, 52)    <= sub_wire17(52);
	sub_wire2(0, 53)    <= sub_wire17(53);
	sub_wire2(0, 54)    <= sub_wire17(54);
	sub_wire2(0, 55)    <= sub_wire17(55);
	sub_wire2(0, 56)    <= sub_wire17(56);
	sub_wire2(0, 57)    <= sub_wire17(57);
	sub_wire2(0, 58)    <= sub_wire17(58);
	sub_wire2(0, 59)    <= sub_wire17(59);
	sub_wire2(0, 60)    <= sub_wire17(60);
	sub_wire2(0, 61)    <= sub_wire17(61);
	sub_wire2(0, 62)    <= sub_wire17(62);
	sub_wire2(0, 63)    <= sub_wire17(63);
	sub_wire2(0, 64)    <= sub_wire17(64);
	sub_wire2(0, 65)    <= sub_wire17(65);
	sub_wire2(0, 66)    <= sub_wire17(66);
	sub_wire2(0, 67)    <= sub_wire17(67);
	sub_wire2(0, 68)    <= sub_wire17(68);
	sub_wire2(0, 69)    <= sub_wire17(69);
	sub_wire2(0, 70)    <= sub_wire17(70);
	sub_wire2(0, 71)    <= sub_wire17(71);
	sub_wire2(0, 72)    <= sub_wire17(72);
	sub_wire2(0, 73)    <= sub_wire17(73);
	sub_wire2(0, 74)    <= sub_wire17(74);
	sub_wire2(0, 75)    <= sub_wire17(75);
	sub_wire2(0, 76)    <= sub_wire17(76);
	sub_wire2(0, 77)    <= sub_wire17(77);
	sub_wire2(0, 78)    <= sub_wire17(78);
	sub_wire2(0, 79)    <= sub_wire17(79);
	sub_wire2(0, 80)    <= sub_wire17(80);
	sub_wire2(0, 81)    <= sub_wire17(81);
	sub_wire2(0, 82)    <= sub_wire17(82);
	sub_wire2(0, 83)    <= sub_wire17(83);
	sub_wire2(0, 84)    <= sub_wire17(84);
	sub_wire2(0, 85)    <= sub_wire17(85);
	sub_wire2(0, 86)    <= sub_wire17(86);
	sub_wire2(0, 87)    <= sub_wire17(87);
	sub_wire2(0, 88)    <= sub_wire17(88);
	sub_wire2(0, 89)    <= sub_wire17(89);
	sub_wire2(0, 90)    <= sub_wire17(90);
	sub_wire2(0, 91)    <= sub_wire17(91);
	sub_wire2(0, 92)    <= sub_wire17(92);
	sub_wire2(0, 93)    <= sub_wire17(93);
	sub_wire2(0, 94)    <= sub_wire17(94);
	sub_wire2(0, 95)    <= sub_wire17(95);
	sub_wire2(0, 96)    <= sub_wire17(96);
	sub_wire2(0, 97)    <= sub_wire17(97);
	sub_wire2(0, 98)    <= sub_wire17(98);
	sub_wire2(0, 99)    <= sub_wire17(99);
	sub_wire2(0, 100)    <= sub_wire17(100);
	sub_wire2(0, 101)    <= sub_wire17(101);
	sub_wire2(0, 102)    <= sub_wire17(102);
	sub_wire2(0, 103)    <= sub_wire17(103);
	sub_wire2(0, 104)    <= sub_wire17(104);
	sub_wire2(0, 105)    <= sub_wire17(105);
	sub_wire2(0, 106)    <= sub_wire17(106);
	sub_wire2(0, 107)    <= sub_wire17(107);
	sub_wire2(0, 108)    <= sub_wire17(108);
	sub_wire2(0, 109)    <= sub_wire17(109);
	sub_wire2(0, 110)    <= sub_wire17(110);
	sub_wire2(0, 111)    <= sub_wire17(111);
	sub_wire2(0, 112)    <= sub_wire17(112);
	sub_wire2(0, 113)    <= sub_wire17(113);
	sub_wire2(0, 114)    <= sub_wire17(114);
	sub_wire2(0, 115)    <= sub_wire17(115);
	sub_wire2(0, 116)    <= sub_wire17(116);
	sub_wire2(0, 117)    <= sub_wire17(117);
	sub_wire2(0, 118)    <= sub_wire17(118);
	sub_wire2(0, 119)    <= sub_wire17(119);
	sub_wire2(0, 120)    <= sub_wire17(120);
	sub_wire2(0, 121)    <= sub_wire17(121);
	sub_wire2(0, 122)    <= sub_wire17(122);
	sub_wire2(0, 123)    <= sub_wire17(123);
	sub_wire2(0, 124)    <= sub_wire17(124);
	sub_wire2(0, 125)    <= sub_wire17(125);
	sub_wire2(0, 126)    <= sub_wire17(126);
	sub_wire2(0, 127)    <= sub_wire17(127);

	lpm_mux_component : lpm_mux
	GENERIC MAP (
		lpm_size => 16,
		lpm_type => "LPM_MUX",
		lpm_width => 128,
		lpm_widths => 4
	)
	PORT MAP (
		sel => sel,
		data => sub_wire2,
		result => sub_wire0
	);



END SYN;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone III"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: CONSTANT: LPM_SIZE NUMERIC "16"
-- Retrieval info: CONSTANT: LPM_TYPE STRING "LPM_MUX"
-- Retrieval info: CONSTANT: LPM_WIDTH NUMERIC "128"
-- Retrieval info: CONSTANT: LPM_WIDTHS NUMERIC "4"
-- Retrieval info: USED_PORT: data0x 0 0 128 0 INPUT NODEFVAL data0x[127..0]
-- Retrieval info: USED_PORT: data10x 0 0 128 0 INPUT NODEFVAL data10x[127..0]
-- Retrieval info: USED_PORT: data11x 0 0 128 0 INPUT NODEFVAL data11x[127..0]
-- Retrieval info: USED_PORT: data12x 0 0 128 0 INPUT NODEFVAL data12x[127..0]
-- Retrieval info: USED_PORT: data13x 0 0 128 0 INPUT NODEFVAL data13x[127..0]
-- Retrieval info: USED_PORT: data14x 0 0 128 0 INPUT NODEFVAL data14x[127..0]
-- Retrieval info: USED_PORT: data15x 0 0 128 0 INPUT NODEFVAL data15x[127..0]
-- Retrieval info: USED_PORT: data1x 0 0 128 0 INPUT NODEFVAL data1x[127..0]
-- Retrieval info: USED_PORT: data2x 0 0 128 0 INPUT NODEFVAL data2x[127..0]
-- Retrieval info: USED_PORT: data3x 0 0 128 0 INPUT NODEFVAL data3x[127..0]
-- Retrieval info: USED_PORT: data4x 0 0 128 0 INPUT NODEFVAL data4x[127..0]
-- Retrieval info: USED_PORT: data5x 0 0 128 0 INPUT NODEFVAL data5x[127..0]
-- Retrieval info: USED_PORT: data6x 0 0 128 0 INPUT NODEFVAL data6x[127..0]
-- Retrieval info: USED_PORT: data7x 0 0 128 0 INPUT NODEFVAL data7x[127..0]
-- Retrieval info: USED_PORT: data8x 0 0 128 0 INPUT NODEFVAL data8x[127..0]
-- Retrieval info: USED_PORT: data9x 0 0 128 0 INPUT NODEFVAL data9x[127..0]
-- Retrieval info: USED_PORT: result 0 0 128 0 OUTPUT NODEFVAL result[127..0]
-- Retrieval info: USED_PORT: sel 0 0 4 0 INPUT NODEFVAL sel[3..0]
-- Retrieval info: CONNECT: result 0 0 128 0 @result 0 0 128 0
-- Retrieval info: CONNECT: @data 1 15 128 0 data15x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 14 128 0 data14x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 13 128 0 data13x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 12 128 0 data12x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 11 128 0 data11x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 10 128 0 data10x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 9 128 0 data9x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 8 128 0 data8x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 7 128 0 data7x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 6 128 0 data6x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 5 128 0 data5x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 4 128 0 data4x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 3 128 0 data3x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 2 128 0 data2x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 1 128 0 data1x 0 0 128 0
-- Retrieval info: CONNECT: @data 1 0 128 0 data0x 0 0 128 0
-- Retrieval info: CONNECT: @sel 0 0 4 0 sel 0 0 4 0
-- Retrieval info: LIBRARY: lpm lpm.lpm_components.all
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_muxVDM.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_muxVDM.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_muxVDM.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_muxVDM.bsf TRUE FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL lpm_muxVDM_inst.vhd FALSE
-- Retrieval info: LIB_FILE: lpm
